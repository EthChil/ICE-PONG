// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Dec 13 2020 21:22:15

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    p_hLED,
    p_vLED,
    p_dwnBtn,
    p_upBtn,
    p_clk12);

    output [14:0] p_hLED;
    output [9:0] p_vLED;
    input p_dwnBtn;
    input p_upBtn;
    input p_clk12;

    wire N__3967;
    wire N__3966;
    wire N__3965;
    wire N__3956;
    wire N__3955;
    wire N__3954;
    wire N__3947;
    wire N__3946;
    wire N__3945;
    wire N__3938;
    wire N__3937;
    wire N__3936;
    wire N__3929;
    wire N__3928;
    wire N__3927;
    wire N__3920;
    wire N__3919;
    wire N__3918;
    wire N__3911;
    wire N__3910;
    wire N__3909;
    wire N__3902;
    wire N__3901;
    wire N__3900;
    wire N__3893;
    wire N__3892;
    wire N__3891;
    wire N__3884;
    wire N__3883;
    wire N__3882;
    wire N__3875;
    wire N__3874;
    wire N__3873;
    wire N__3866;
    wire N__3865;
    wire N__3864;
    wire N__3857;
    wire N__3856;
    wire N__3855;
    wire N__3848;
    wire N__3847;
    wire N__3846;
    wire N__3839;
    wire N__3838;
    wire N__3837;
    wire N__3830;
    wire N__3829;
    wire N__3828;
    wire N__3821;
    wire N__3820;
    wire N__3819;
    wire N__3812;
    wire N__3811;
    wire N__3810;
    wire N__3803;
    wire N__3802;
    wire N__3801;
    wire N__3794;
    wire N__3793;
    wire N__3792;
    wire N__3785;
    wire N__3784;
    wire N__3783;
    wire N__3776;
    wire N__3775;
    wire N__3774;
    wire N__3767;
    wire N__3766;
    wire N__3765;
    wire N__3758;
    wire N__3757;
    wire N__3756;
    wire N__3749;
    wire N__3748;
    wire N__3747;
    wire N__3740;
    wire N__3739;
    wire N__3738;
    wire N__3721;
    wire N__3718;
    wire N__3715;
    wire N__3712;
    wire N__3709;
    wire N__3706;
    wire N__3703;
    wire N__3700;
    wire N__3697;
    wire N__3694;
    wire N__3691;
    wire N__3688;
    wire N__3685;
    wire N__3682;
    wire N__3679;
    wire N__3676;
    wire N__3673;
    wire N__3670;
    wire N__3667;
    wire N__3664;
    wire N__3661;
    wire N__3658;
    wire N__3655;
    wire N__3652;
    wire N__3649;
    wire N__3646;
    wire N__3643;
    wire N__3640;
    wire N__3637;
    wire N__3634;
    wire N__3631;
    wire N__3628;
    wire N__3625;
    wire N__3622;
    wire N__3619;
    wire N__3616;
    wire N__3613;
    wire N__3610;
    wire N__3607;
    wire N__3604;
    wire N__3601;
    wire N__3598;
    wire N__3595;
    wire N__3592;
    wire N__3589;
    wire N__3586;
    wire N__3585;
    wire N__3584;
    wire N__3583;
    wire N__3582;
    wire N__3581;
    wire N__3580;
    wire N__3577;
    wire N__3576;
    wire N__3575;
    wire N__3574;
    wire N__3573;
    wire N__3572;
    wire N__3571;
    wire N__3570;
    wire N__3569;
    wire N__3568;
    wire N__3567;
    wire N__3566;
    wire N__3565;
    wire N__3564;
    wire N__3563;
    wire N__3550;
    wire N__3547;
    wire N__3538;
    wire N__3535;
    wire N__3526;
    wire N__3515;
    wire N__3512;
    wire N__3509;
    wire N__3504;
    wire N__3493;
    wire N__3492;
    wire N__3491;
    wire N__3490;
    wire N__3489;
    wire N__3488;
    wire N__3487;
    wire N__3486;
    wire N__3485;
    wire N__3484;
    wire N__3483;
    wire N__3482;
    wire N__3481;
    wire N__3480;
    wire N__3467;
    wire N__3458;
    wire N__3457;
    wire N__3456;
    wire N__3455;
    wire N__3452;
    wire N__3451;
    wire N__3444;
    wire N__3441;
    wire N__3438;
    wire N__3431;
    wire N__3428;
    wire N__3425;
    wire N__3412;
    wire N__3411;
    wire N__3410;
    wire N__3409;
    wire N__3408;
    wire N__3407;
    wire N__3406;
    wire N__3405;
    wire N__3404;
    wire N__3403;
    wire N__3402;
    wire N__3401;
    wire N__3400;
    wire N__3399;
    wire N__3396;
    wire N__3393;
    wire N__3390;
    wire N__3387;
    wire N__3384;
    wire N__3381;
    wire N__3380;
    wire N__3379;
    wire N__3376;
    wire N__3373;
    wire N__3370;
    wire N__3367;
    wire N__3364;
    wire N__3351;
    wire N__3342;
    wire N__3341;
    wire N__3338;
    wire N__3337;
    wire N__3334;
    wire N__3329;
    wire N__3324;
    wire N__3321;
    wire N__3318;
    wire N__3315;
    wire N__3312;
    wire N__3309;
    wire N__3292;
    wire N__3291;
    wire N__3290;
    wire N__3289;
    wire N__3286;
    wire N__3285;
    wire N__3284;
    wire N__3283;
    wire N__3282;
    wire N__3281;
    wire N__3280;
    wire N__3277;
    wire N__3274;
    wire N__3271;
    wire N__3262;
    wire N__3249;
    wire N__3248;
    wire N__3247;
    wire N__3246;
    wire N__3245;
    wire N__3244;
    wire N__3243;
    wire N__3242;
    wire N__3241;
    wire N__3240;
    wire N__3239;
    wire N__3234;
    wire N__3231;
    wire N__3230;
    wire N__3225;
    wire N__3220;
    wire N__3213;
    wire N__3210;
    wire N__3207;
    wire N__3204;
    wire N__3201;
    wire N__3198;
    wire N__3181;
    wire N__3180;
    wire N__3179;
    wire N__3178;
    wire N__3177;
    wire N__3176;
    wire N__3175;
    wire N__3174;
    wire N__3173;
    wire N__3172;
    wire N__3171;
    wire N__3170;
    wire N__3169;
    wire N__3142;
    wire N__3139;
    wire N__3136;
    wire N__3135;
    wire N__3132;
    wire N__3131;
    wire N__3128;
    wire N__3125;
    wire N__3122;
    wire N__3119;
    wire N__3114;
    wire N__3109;
    wire N__3106;
    wire N__3103;
    wire N__3100;
    wire N__3097;
    wire N__3094;
    wire N__3091;
    wire N__3088;
    wire N__3085;
    wire N__3082;
    wire N__3079;
    wire N__3076;
    wire N__3073;
    wire N__3072;
    wire N__3071;
    wire N__3070;
    wire N__3067;
    wire N__3064;
    wire N__3063;
    wire N__3062;
    wire N__3059;
    wire N__3056;
    wire N__3051;
    wire N__3048;
    wire N__3045;
    wire N__3038;
    wire N__3035;
    wire N__3032;
    wire N__3031;
    wire N__3030;
    wire N__3029;
    wire N__3028;
    wire N__3025;
    wire N__3020;
    wire N__3017;
    wire N__3014;
    wire N__3011;
    wire N__3008;
    wire N__2995;
    wire N__2992;
    wire N__2989;
    wire N__2986;
    wire N__2983;
    wire N__2980;
    wire N__2977;
    wire N__2974;
    wire N__2973;
    wire N__2972;
    wire N__2967;
    wire N__2964;
    wire N__2959;
    wire N__2956;
    wire N__2953;
    wire N__2950;
    wire N__2947;
    wire N__2944;
    wire N__2941;
    wire N__2938;
    wire N__2935;
    wire N__2932;
    wire N__2929;
    wire N__2926;
    wire N__2923;
    wire N__2920;
    wire N__2917;
    wire N__2914;
    wire N__2911;
    wire N__2908;
    wire N__2905;
    wire N__2902;
    wire N__2899;
    wire N__2896;
    wire N__2893;
    wire N__2890;
    wire N__2887;
    wire N__2884;
    wire N__2881;
    wire N__2878;
    wire N__2875;
    wire N__2872;
    wire N__2869;
    wire N__2866;
    wire N__2863;
    wire N__2860;
    wire N__2857;
    wire N__2854;
    wire N__2851;
    wire N__2848;
    wire N__2845;
    wire N__2842;
    wire N__2839;
    wire N__2836;
    wire N__2833;
    wire N__2830;
    wire N__2827;
    wire N__2824;
    wire N__2821;
    wire N__2818;
    wire N__2815;
    wire N__2812;
    wire N__2811;
    wire N__2810;
    wire N__2807;
    wire N__2804;
    wire N__2801;
    wire N__2798;
    wire N__2791;
    wire N__2790;
    wire N__2787;
    wire N__2786;
    wire N__2783;
    wire N__2780;
    wire N__2777;
    wire N__2774;
    wire N__2771;
    wire N__2764;
    wire N__2763;
    wire N__2762;
    wire N__2759;
    wire N__2754;
    wire N__2751;
    wire N__2746;
    wire N__2743;
    wire N__2740;
    wire N__2737;
    wire N__2734;
    wire N__2731;
    wire N__2728;
    wire N__2727;
    wire N__2726;
    wire N__2723;
    wire N__2718;
    wire N__2715;
    wire N__2710;
    wire N__2709;
    wire N__2706;
    wire N__2703;
    wire N__2700;
    wire N__2695;
    wire N__2692;
    wire N__2689;
    wire N__2688;
    wire N__2685;
    wire N__2682;
    wire N__2679;
    wire N__2674;
    wire N__2671;
    wire N__2668;
    wire N__2667;
    wire N__2664;
    wire N__2661;
    wire N__2658;
    wire N__2653;
    wire N__2650;
    wire N__2647;
    wire N__2646;
    wire N__2643;
    wire N__2640;
    wire N__2637;
    wire N__2632;
    wire N__2629;
    wire N__2626;
    wire N__2623;
    wire N__2620;
    wire N__2617;
    wire N__2614;
    wire N__2611;
    wire N__2608;
    wire N__2605;
    wire N__2602;
    wire N__2599;
    wire N__2596;
    wire N__2593;
    wire N__2590;
    wire N__2587;
    wire N__2584;
    wire N__2581;
    wire N__2578;
    wire N__2575;
    wire N__2572;
    wire N__2569;
    wire N__2566;
    wire N__2563;
    wire N__2560;
    wire N__2557;
    wire N__2554;
    wire N__2551;
    wire N__2548;
    wire N__2545;
    wire N__2542;
    wire N__2539;
    wire N__2538;
    wire N__2535;
    wire N__2532;
    wire N__2529;
    wire N__2524;
    wire N__2521;
    wire N__2518;
    wire N__2517;
    wire N__2514;
    wire N__2511;
    wire N__2506;
    wire N__2503;
    wire N__2502;
    wire N__2499;
    wire N__2496;
    wire N__2493;
    wire N__2488;
    wire N__2485;
    wire N__2484;
    wire N__2481;
    wire N__2478;
    wire N__2473;
    wire N__2470;
    wire N__2469;
    wire N__2466;
    wire N__2463;
    wire N__2458;
    wire N__2455;
    wire N__2454;
    wire N__2451;
    wire N__2448;
    wire N__2443;
    wire N__2440;
    wire N__2439;
    wire N__2436;
    wire N__2433;
    wire N__2428;
    wire N__2425;
    wire N__2424;
    wire N__2421;
    wire N__2418;
    wire N__2415;
    wire N__2410;
    wire N__2407;
    wire N__2406;
    wire N__2405;
    wire N__2404;
    wire N__2401;
    wire N__2398;
    wire N__2395;
    wire N__2392;
    wire N__2383;
    wire N__2380;
    wire N__2377;
    wire N__2376;
    wire N__2373;
    wire N__2370;
    wire N__2365;
    wire N__2364;
    wire N__2363;
    wire N__2362;
    wire N__2361;
    wire N__2360;
    wire N__2359;
    wire N__2346;
    wire N__2345;
    wire N__2344;
    wire N__2343;
    wire N__2340;
    wire N__2339;
    wire N__2338;
    wire N__2335;
    wire N__2328;
    wire N__2325;
    wire N__2320;
    wire N__2311;
    wire N__2310;
    wire N__2307;
    wire N__2304;
    wire N__2299;
    wire N__2296;
    wire N__2293;
    wire N__2292;
    wire N__2289;
    wire N__2286;
    wire N__2283;
    wire N__2278;
    wire N__2275;
    wire N__2274;
    wire N__2271;
    wire N__2268;
    wire N__2263;
    wire N__2260;
    wire N__2259;
    wire N__2256;
    wire N__2253;
    wire N__2248;
    wire N__2245;
    wire N__2244;
    wire N__2241;
    wire N__2238;
    wire N__2233;
    wire N__2230;
    wire N__2229;
    wire N__2226;
    wire N__2223;
    wire N__2218;
    wire N__2215;
    wire N__2214;
    wire N__2211;
    wire N__2208;
    wire N__2205;
    wire N__2200;
    wire N__2197;
    wire N__2194;
    wire N__2191;
    wire N__2188;
    wire N__2185;
    wire N__2182;
    wire N__2179;
    wire N__2178;
    wire N__2175;
    wire N__2172;
    wire N__2169;
    wire N__2166;
    wire N__2161;
    wire N__2160;
    wire N__2159;
    wire N__2158;
    wire N__2157;
    wire N__2156;
    wire N__2155;
    wire N__2154;
    wire N__2141;
    wire N__2140;
    wire N__2139;
    wire N__2138;
    wire N__2135;
    wire N__2134;
    wire N__2131;
    wire N__2128;
    wire N__2121;
    wire N__2116;
    wire N__2113;
    wire N__2104;
    wire N__2103;
    wire N__2102;
    wire N__2101;
    wire N__2100;
    wire N__2097;
    wire N__2094;
    wire N__2091;
    wire N__2090;
    wire N__2089;
    wire N__2088;
    wire N__2085;
    wire N__2082;
    wire N__2081;
    wire N__2068;
    wire N__2067;
    wire N__2066;
    wire N__2065;
    wire N__2058;
    wire N__2055;
    wire N__2052;
    wire N__2049;
    wire N__2046;
    wire N__2035;
    wire N__2034;
    wire N__2033;
    wire N__2032;
    wire N__2031;
    wire N__2030;
    wire N__2027;
    wire N__2024;
    wire N__2021;
    wire N__2020;
    wire N__2019;
    wire N__2006;
    wire N__2005;
    wire N__2004;
    wire N__2001;
    wire N__2000;
    wire N__1999;
    wire N__1996;
    wire N__1993;
    wire N__1986;
    wire N__1983;
    wire N__1980;
    wire N__1977;
    wire N__1966;
    wire N__1963;
    wire N__1960;
    wire N__1957;
    wire N__1954;
    wire N__1951;
    wire N__1948;
    wire N__1945;
    wire N__1942;
    wire N__1939;
    wire N__1938;
    wire N__1937;
    wire N__1936;
    wire N__1933;
    wire N__1932;
    wire N__1931;
    wire N__1928;
    wire N__1927;
    wire N__1926;
    wire N__1925;
    wire N__1922;
    wire N__1921;
    wire N__1918;
    wire N__1913;
    wire N__1904;
    wire N__1897;
    wire N__1888;
    wire N__1885;
    wire N__1882;
    wire N__1879;
    wire N__1876;
    wire N__1873;
    wire N__1870;
    wire N__1867;
    wire N__1864;
    wire N__1861;
    wire N__1858;
    wire N__1855;
    wire N__1852;
    wire N__1849;
    wire N__1848;
    wire N__1847;
    wire N__1844;
    wire N__1839;
    wire N__1834;
    wire N__1831;
    wire N__1830;
    wire N__1829;
    wire N__1826;
    wire N__1823;
    wire N__1820;
    wire N__1813;
    wire N__1810;
    wire N__1809;
    wire N__1808;
    wire N__1807;
    wire N__1806;
    wire N__1803;
    wire N__1798;
    wire N__1793;
    wire N__1786;
    wire N__1785;
    wire N__1782;
    wire N__1781;
    wire N__1778;
    wire N__1773;
    wire N__1768;
    wire N__1767;
    wire N__1764;
    wire N__1763;
    wire N__1760;
    wire N__1757;
    wire N__1752;
    wire N__1747;
    wire N__1744;
    wire N__1741;
    wire N__1738;
    wire N__1735;
    wire N__1732;
    wire N__1729;
    wire N__1726;
    wire N__1723;
    wire N__1720;
    wire N__1717;
    wire N__1716;
    wire N__1715;
    wire N__1714;
    wire N__1713;
    wire N__1702;
    wire N__1699;
    wire N__1696;
    wire N__1693;
    wire N__1690;
    wire N__1687;
    wire N__1684;
    wire N__1681;
    wire N__1678;
    wire N__1675;
    wire N__1672;
    wire N__1669;
    wire N__1666;
    wire VCCG0;
    wire GNDG0;
    wire bfn_7_6_0_;
    wire un1_ballY_4_cry_0;
    wire un1_ballY_4_cry_1;
    wire un1_ballY_4_cry_2;
    wire ballYVel_RNIGOGN4_0Z0Z_0;
    wire ballYVel_RNIGOGN4Z0Z_0;
    wire bfn_7_7_0_;
    wire un1_ballX_3_cry_0;
    wire un1_ballX_3_cry_1;
    wire un1_ballX_3_cry_2;
    wire ballXVel_s_1_0_0_cascade_;
    wire ballXVel_RNIFI1J4_0Z0Z_0;
    wire ballXVelZ0Z_0;
    wire ballXVel_RNIFI1J4Z0Z_0;
    wire N_67_i;
    wire bfn_8_6_0_;
    wire un1_vIndex_2_cry_0;
    wire un1_vIndex_2_cry_1;
    wire un1_vIndex_2_cry_2;
    wire ballYZ0Z_0;
    wire ballYZ0Z_1;
    wire ballYVel_s_1_0_0_cascade_;
    wire ballYVelZ0Z_0;
    wire ballYZ0Z_2;
    wire ballYZ0Z_3;
    wire p_vLED37_NE_0;
    wire ballXVel12_10_cascade_;
    wire ballXVel12_12;
    wire ballXVel12_14_cascade_;
    wire ballXVel12_11;
    wire ballXVel12;
    wire ballXVel12_13;
    wire N_430_i;
    wire N_428_i;
    wire p_vLED_cl_2_iZ0Z_0;
    wire p_vLED_cl_9_iZ0Z_0;
    wire p_vLED37;
    wire vIndexZ0Z_2;
    wire vIndexZ0Z_1;
    wire vIndexZ0Z_3;
    wire N_76_cascade_;
    wire N_57_i;
    wire p_vLED33;
    wire N_57_i_cascade_;
    wire N_76;
    wire vIndexZ0Z_0;
    wire ctrZ0Z_0;
    wire bfn_9_7_0_;
    wire ctrZ0Z_1;
    wire ctr_cry_0;
    wire ctrZ0Z_2;
    wire ctr_cry_1;
    wire ctrZ0Z_3;
    wire ctr_cry_2;
    wire ctrZ0Z_4;
    wire ctr_cry_3;
    wire ctrZ0Z_5;
    wire ctr_cry_4;
    wire ctrZ0Z_6;
    wire ctr_cry_5;
    wire ctrZ0Z_7;
    wire ctr_cry_6;
    wire ctr_cry_7;
    wire ctrZ0Z_8;
    wire bfn_9_8_0_;
    wire ctrZ0Z_9;
    wire ctr_cry_8;
    wire ctrZ0Z_10;
    wire ctr_cry_9;
    wire ctrZ0Z_11;
    wire ctr_cry_10;
    wire ctrZ0Z_12;
    wire ctr_cry_11;
    wire ctrZ0Z_13;
    wire ctr_cry_12;
    wire ctrZ0Z_14;
    wire ctr_cry_13;
    wire ctrZ0Z_15;
    wire ctr_cry_14;
    wire ctr_cry_15;
    wire ctrZ0Z_16;
    wire bfn_9_9_0_;
    wire ctrZ0Z_17;
    wire ctr_cry_16;
    wire ctr_cry_17;
    wire ctrZ0Z_18;
    wire N_412_i;
    wire p_vLED_cl_iZ0Z_0;
    wire N_429_i;
    wire p_vLED_cl_6_iZ0Z_0;
    wire N_425_i;
    wire p_vLED_cl_8_iZ0Z_0;
    wire N_424_i;
    wire p_vLED_cl_3_iZ0Z_0;
    wire N_422_i;
    wire N_58_cascade_;
    wire p_vLED_cl_1_iZ0Z_0;
    wire N_423_i;
    wire ballXZ0Z_1;
    wire ballXZ0Z_2;
    wire ballXZ0Z_0;
    wire p_hLED52_NE_0;
    wire N_70_i;
    wire ballXZ0Z_3;
    wire N_410_i;
    wire p_hLED_cl_6_iZ0Z_0;
    wire p_vLED_cl_4_iZ0Z_0;
    wire N_427_i;
    wire p_vLED_cl_7_iZ0Z_0;
    wire N_426_i;
    wire N_414_i;
    wire p_vLED_cl_5_iZ0Z_0;
    wire N_421_i;
    wire CONSTANT_ONE_NET;
    wire p_hLED_cl_7_iZ0Z_0;
    wire p_hLED_cl_iZ0Z_0;
    wire N_58;
    wire p_hLED_cl_14_iZ0Z_0;
    wire N_406_i;
    wire p_hLED_cl_4_iZ0Z_0;
    wire N_408_i;
    wire N_407_i;
    wire p_hLED_cl_2_iZ0Z_0;
    wire N_409_i;
    wire p_hLED_cl_3_iZ0Z_0;
    wire hIndexZ0Z_3;
    wire hIndexZ0Z_2;
    wire hIndexZ0Z_1;
    wire hIndexZ0Z_0;
    wire p_clk12_c_g;
    wire p_hLED52;
    wire p_hLED_cl_13_iZ0Z_0;
    wire N_416_i;
    wire p_hLED_cl_8_iZ0Z_0;
    wire N_411_i;
    wire p_hLED_cl_10_iZ0Z_0;
    wire N_417_i;
    wire p_hLED_cl_9_iZ0Z_0;
    wire N_418_i;
    wire p_hLED_cl_1_iZ0Z_0;
    wire N_413_i;
    wire p_hLED_cl_11_iZ0Z_0;
    wire N_420_i;
    wire p_hLED_cl_12_iZ0Z_0;
    wire N_415_i;
    wire p_hLED_cl_5_iZ0Z_0;
    wire N_419_i;
    wire _gnd_net_;

    PRE_IO_GBUF p_clk12_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__3965),
            .GLOBALBUFFEROUTPUT(p_clk12_c_g));
    defparam p_clk12_ibuf_gb_io_iopad.PULLUP=1'b0;
    defparam p_clk12_ibuf_gb_io_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD p_clk12_ibuf_gb_io_iopad (
            .OE(N__3967),
            .DIN(N__3966),
            .DOUT(N__3965),
            .PACKAGEPIN(p_clk12));
    defparam p_clk12_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam p_clk12_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO p_clk12_ibuf_gb_io_preio (
            .PADOEN(N__3967),
            .PADOUT(N__3966),
            .PADIN(N__3965),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam p_vLED_obuft_0_iopad.PULLUP=1'b0;
    defparam p_vLED_obuft_0_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD p_vLED_obuft_0_iopad (
            .OE(N__3956),
            .DIN(N__3955),
            .DOUT(N__3954),
            .PACKAGEPIN(p_vLED[0]));
    defparam p_vLED_obuft_0_preio.NEG_TRIGGER=1'b0;
    defparam p_vLED_obuft_0_preio.PIN_TYPE=6'b101001;
    PRE_IO p_vLED_obuft_0_preio (
            .PADOEN(N__3956),
            .PADOUT(N__3955),
            .PADIN(N__3954),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2851),
            .DIN0(),
            .DOUT0(N__3063),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam p_hLED_obuft_2_iopad.PULLUP=1'b0;
    defparam p_hLED_obuft_2_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD p_hLED_obuft_2_iopad (
            .OE(N__3947),
            .DIN(N__3946),
            .DOUT(N__3945),
            .PACKAGEPIN(p_hLED[2]));
    defparam p_hLED_obuft_2_preio.NEG_TRIGGER=1'b0;
    defparam p_hLED_obuft_2_preio.PIN_TYPE=6'b101001;
    PRE_IO p_hLED_obuft_2_preio (
            .PADOEN(N__3947),
            .PADOUT(N__3946),
            .PADIN(N__3945),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2941),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam p_hLED_obuft_5_iopad.PULLUP=1'b0;
    defparam p_hLED_obuft_5_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD p_hLED_obuft_5_iopad (
            .OE(N__3938),
            .DIN(N__3937),
            .DOUT(N__3936),
            .PACKAGEPIN(p_hLED[5]));
    defparam p_hLED_obuft_5_preio.NEG_TRIGGER=1'b0;
    defparam p_hLED_obuft_5_preio.PIN_TYPE=6'b101001;
    PRE_IO p_hLED_obuft_5_preio (
            .PADOEN(N__3938),
            .PADOUT(N__3937),
            .PADIN(N__3936),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3079),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam p_hLED_obuft_10_iopad.PULLUP=1'b0;
    defparam p_hLED_obuft_10_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD p_hLED_obuft_10_iopad (
            .OE(N__3929),
            .DIN(N__3928),
            .DOUT(N__3927),
            .PACKAGEPIN(p_hLED[10]));
    defparam p_hLED_obuft_10_preio.NEG_TRIGGER=1'b0;
    defparam p_hLED_obuft_10_preio.PIN_TYPE=6'b101001;
    PRE_IO p_hLED_obuft_10_preio (
            .PADOEN(N__3929),
            .PADOUT(N__3928),
            .PADIN(N__3927),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3097),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam p_vLED_obuft_7_iopad.PULLUP=1'b0;
    defparam p_vLED_obuft_7_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD p_vLED_obuft_7_iopad (
            .OE(N__3920),
            .DIN(N__3919),
            .DOUT(N__3918),
            .PACKAGEPIN(p_vLED[7]));
    defparam p_vLED_obuft_7_preio.NEG_TRIGGER=1'b0;
    defparam p_vLED_obuft_7_preio.PIN_TYPE=6'b101001;
    PRE_IO p_vLED_obuft_7_preio (
            .PADOEN(N__3920),
            .PADOUT(N__3919),
            .PADIN(N__3918),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__1873),
            .DIN0(),
            .DOUT0(N__3072),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam p_vLED_obuft_2_iopad.PULLUP=1'b0;
    defparam p_vLED_obuft_2_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD p_vLED_obuft_2_iopad (
            .OE(N__3911),
            .DIN(N__3910),
            .DOUT(N__3909),
            .PACKAGEPIN(p_vLED[2]));
    defparam p_vLED_obuft_2_preio.NEG_TRIGGER=1'b0;
    defparam p_vLED_obuft_2_preio.PIN_TYPE=6'b101001;
    PRE_IO p_vLED_obuft_2_preio (
            .PADOEN(N__3911),
            .PADOUT(N__3910),
            .PADIN(N__3909),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2821),
            .DIN0(),
            .DOUT0(N__3030),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam p_vLED_obuft_9_iopad.PULLUP=1'b0;
    defparam p_vLED_obuft_9_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD p_vLED_obuft_9_iopad (
            .OE(N__3902),
            .DIN(N__3901),
            .DOUT(N__3900),
            .PACKAGEPIN(p_vLED[9]));
    defparam p_vLED_obuft_9_preio.NEG_TRIGGER=1'b0;
    defparam p_vLED_obuft_9_preio.PIN_TYPE=6'b101001;
    PRE_IO p_vLED_obuft_9_preio (
            .PADOEN(N__3902),
            .PADOUT(N__3901),
            .PADIN(N__3900),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__1882),
            .DIN0(),
            .DOUT0(N__3070),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam p_hLED_obuft_0_iopad.PULLUP=1'b0;
    defparam p_hLED_obuft_0_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD p_hLED_obuft_0_iopad (
            .OE(N__3893),
            .DIN(N__3892),
            .DOUT(N__3891),
            .PACKAGEPIN(p_hLED[0]));
    defparam p_hLED_obuft_0_preio.NEG_TRIGGER=1'b0;
    defparam p_hLED_obuft_0_preio.PIN_TYPE=6'b101001;
    PRE_IO p_hLED_obuft_0_preio (
            .PADOEN(N__3893),
            .PADOUT(N__3892),
            .PADIN(N__3891),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2953),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam p_vLED_obuft_1_iopad.PULLUP=1'b0;
    defparam p_vLED_obuft_1_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD p_vLED_obuft_1_iopad (
            .OE(N__3884),
            .DIN(N__3883),
            .DOUT(N__3882),
            .PACKAGEPIN(p_vLED[1]));
    defparam p_vLED_obuft_1_preio.NEG_TRIGGER=1'b0;
    defparam p_vLED_obuft_1_preio.PIN_TYPE=6'b101001;
    PRE_IO p_vLED_obuft_1_preio (
            .PADOEN(N__3884),
            .PADOUT(N__3883),
            .PADIN(N__3882),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2551),
            .DIN0(),
            .DOUT0(N__3031),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam p_hLED_obuft_7_iopad.PULLUP=1'b0;
    defparam p_hLED_obuft_7_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD p_hLED_obuft_7_iopad (
            .OE(N__3875),
            .DIN(N__3874),
            .DOUT(N__3873),
            .PACKAGEPIN(p_hLED[7]));
    defparam p_hLED_obuft_7_preio.NEG_TRIGGER=1'b0;
    defparam p_hLED_obuft_7_preio.PIN_TYPE=6'b101001;
    PRE_IO p_hLED_obuft_7_preio (
            .PADOEN(N__3875),
            .PADOUT(N__3874),
            .PADIN(N__3873),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3664),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam p_hLED_obuft_12_iopad.PULLUP=1'b0;
    defparam p_hLED_obuft_12_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD p_hLED_obuft_12_iopad (
            .OE(N__3866),
            .DIN(N__3865),
            .DOUT(N__3864),
            .PACKAGEPIN(p_hLED[12]));
    defparam p_hLED_obuft_12_preio.NEG_TRIGGER=1'b0;
    defparam p_hLED_obuft_12_preio.PIN_TYPE=6'b101001;
    PRE_IO p_hLED_obuft_12_preio (
            .PADOEN(N__3866),
            .PADOUT(N__3865),
            .PADIN(N__3864),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3691),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam p_hLED_obuft_8_iopad.PULLUP=1'b0;
    defparam p_hLED_obuft_8_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD p_hLED_obuft_8_iopad (
            .OE(N__3857),
            .DIN(N__3856),
            .DOUT(N__3855),
            .PACKAGEPIN(p_hLED[8]));
    defparam p_hLED_obuft_8_preio.NEG_TRIGGER=1'b0;
    defparam p_hLED_obuft_8_preio.PIN_TYPE=6'b101001;
    PRE_IO p_hLED_obuft_8_preio (
            .PADOEN(N__3857),
            .PADOUT(N__3856),
            .PADIN(N__3855),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2872),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam p_vLED_obuft_5_iopad.PULLUP=1'b0;
    defparam p_vLED_obuft_5_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD p_vLED_obuft_5_iopad (
            .OE(N__3848),
            .DIN(N__3847),
            .DOUT(N__3846),
            .PACKAGEPIN(p_vLED[5]));
    defparam p_vLED_obuft_5_preio.NEG_TRIGGER=1'b0;
    defparam p_vLED_obuft_5_preio.PIN_TYPE=6'b101001;
    PRE_IO p_vLED_obuft_5_preio (
            .PADOEN(N__3848),
            .PADOUT(N__3847),
            .PADIN(N__3846),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2878),
            .DIN0(),
            .DOUT0(N__3062),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam p_hLED_obuft_3_iopad.PULLUP=1'b0;
    defparam p_hLED_obuft_3_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD p_hLED_obuft_3_iopad (
            .OE(N__3839),
            .DIN(N__3838),
            .DOUT(N__3837),
            .PACKAGEPIN(p_hLED[3]));
    defparam p_hLED_obuft_3_preio.NEG_TRIGGER=1'b0;
    defparam p_hLED_obuft_3_preio.PIN_TYPE=6'b101001;
    PRE_IO p_hLED_obuft_3_preio (
            .PADOEN(N__3839),
            .PADOUT(N__3838),
            .PADIN(N__3837),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3598),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam p_hLED_obuft_6_iopad.PULLUP=1'b0;
    defparam p_hLED_obuft_6_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD p_hLED_obuft_6_iopad (
            .OE(N__3830),
            .DIN(N__3829),
            .DOUT(N__3828),
            .PACKAGEPIN(p_hLED[6]));
    defparam p_hLED_obuft_6_preio.NEG_TRIGGER=1'b0;
    defparam p_hLED_obuft_6_preio.PIN_TYPE=6'b101001;
    PRE_IO p_hLED_obuft_6_preio (
            .PADOEN(N__3830),
            .PADOUT(N__3829),
            .PADIN(N__3828),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2632),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam p_hLED_obuft_13_iopad.PULLUP=1'b0;
    defparam p_hLED_obuft_13_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD p_hLED_obuft_13_iopad (
            .OE(N__3821),
            .DIN(N__3820),
            .DOUT(N__3819),
            .PACKAGEPIN(p_hLED[13]));
    defparam p_hLED_obuft_13_preio.NEG_TRIGGER=1'b0;
    defparam p_hLED_obuft_13_preio.PIN_TYPE=6'b101001;
    PRE_IO p_hLED_obuft_13_preio (
            .PADOEN(N__3821),
            .PADOUT(N__3820),
            .PADIN(N__3819),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3610),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam p_vLED_obuft_4_iopad.PULLUP=1'b0;
    defparam p_vLED_obuft_4_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD p_vLED_obuft_4_iopad (
            .OE(N__3812),
            .DIN(N__3811),
            .DOUT(N__3810),
            .PACKAGEPIN(p_vLED[4]));
    defparam p_vLED_obuft_4_preio.NEG_TRIGGER=1'b0;
    defparam p_vLED_obuft_4_preio.PIN_TYPE=6'b101001;
    PRE_IO p_vLED_obuft_4_preio (
            .PADOEN(N__3812),
            .PADOUT(N__3811),
            .PADIN(N__3810),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2587),
            .DIN0(),
            .DOUT0(N__3028),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam p_vLED_obuft_3_iopad.PULLUP=1'b0;
    defparam p_vLED_obuft_3_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD p_vLED_obuft_3_iopad (
            .OE(N__3803),
            .DIN(N__3802),
            .DOUT(N__3801),
            .PACKAGEPIN(p_vLED[3]));
    defparam p_vLED_obuft_3_preio.NEG_TRIGGER=1'b0;
    defparam p_vLED_obuft_3_preio.PIN_TYPE=6'b101001;
    PRE_IO p_vLED_obuft_3_preio (
            .PADOEN(N__3803),
            .PADOUT(N__3802),
            .PADIN(N__3801),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2569),
            .DIN0(),
            .DOUT0(N__3029),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam p_hLED_obuft_1_iopad.PULLUP=1'b0;
    defparam p_hLED_obuft_1_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD p_hLED_obuft_1_iopad (
            .OE(N__3794),
            .DIN(N__3793),
            .DOUT(N__3792),
            .PACKAGEPIN(p_hLED[1]));
    defparam p_hLED_obuft_1_preio.NEG_TRIGGER=1'b0;
    defparam p_hLED_obuft_1_preio.PIN_TYPE=6'b101001;
    PRE_IO p_hLED_obuft_1_preio (
            .PADOEN(N__3794),
            .PADOUT(N__3793),
            .PADIN(N__3792),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2935),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam p_hLED_obuft_14_iopad.PULLUP=1'b0;
    defparam p_hLED_obuft_14_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD p_hLED_obuft_14_iopad (
            .OE(N__3785),
            .DIN(N__3784),
            .DOUT(N__3783),
            .PACKAGEPIN(p_hLED[14]));
    defparam p_hLED_obuft_14_preio.NEG_TRIGGER=1'b0;
    defparam p_hLED_obuft_14_preio.PIN_TYPE=6'b101001;
    PRE_IO p_hLED_obuft_14_preio (
            .PADOEN(N__3785),
            .PADOUT(N__3784),
            .PADIN(N__3783),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3649),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam p_hLED_obuft_4_iopad.PULLUP=1'b0;
    defparam p_hLED_obuft_4_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD p_hLED_obuft_4_iopad (
            .OE(N__3776),
            .DIN(N__3775),
            .DOUT(N__3774),
            .PACKAGEPIN(p_hLED[4]));
    defparam p_hLED_obuft_4_preio.NEG_TRIGGER=1'b0;
    defparam p_hLED_obuft_4_preio.PIN_TYPE=6'b101001;
    PRE_IO p_hLED_obuft_4_preio (
            .PADOEN(N__3776),
            .PADOUT(N__3775),
            .PADIN(N__3774),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2929),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam p_hLED_obuft_11_iopad.PULLUP=1'b0;
    defparam p_hLED_obuft_11_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD p_hLED_obuft_11_iopad (
            .OE(N__3767),
            .DIN(N__3766),
            .DOUT(N__3765),
            .PACKAGEPIN(p_hLED[11]));
    defparam p_hLED_obuft_11_preio.NEG_TRIGGER=1'b0;
    defparam p_hLED_obuft_11_preio.PIN_TYPE=6'b101001;
    PRE_IO p_hLED_obuft_11_preio (
            .PADOEN(N__3767),
            .PADOUT(N__3766),
            .PADIN(N__3765),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3715),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam p_vLED_obuft_6_iopad.PULLUP=1'b0;
    defparam p_vLED_obuft_6_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD p_vLED_obuft_6_iopad (
            .OE(N__3758),
            .DIN(N__3757),
            .DOUT(N__3756),
            .PACKAGEPIN(p_vLED[6]));
    defparam p_vLED_obuft_6_preio.NEG_TRIGGER=1'b0;
    defparam p_vLED_obuft_6_preio.PIN_TYPE=6'b101001;
    PRE_IO p_vLED_obuft_6_preio (
            .PADOEN(N__3758),
            .PADOUT(N__3757),
            .PADIN(N__3756),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2896),
            .DIN0(),
            .DOUT0(N__3073),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam p_hLED_obuft_9_iopad.PULLUP=1'b0;
    defparam p_hLED_obuft_9_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD p_hLED_obuft_9_iopad (
            .OE(N__3749),
            .DIN(N__3748),
            .DOUT(N__3747),
            .PACKAGEPIN(p_hLED[9]));
    defparam p_hLED_obuft_9_preio.NEG_TRIGGER=1'b0;
    defparam p_hLED_obuft_9_preio.PIN_TYPE=6'b101001;
    PRE_IO p_hLED_obuft_9_preio (
            .PADOEN(N__3749),
            .PADOUT(N__3748),
            .PADIN(N__3747),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3625),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam p_vLED_obuft_8_iopad.PULLUP=1'b0;
    defparam p_vLED_obuft_8_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD p_vLED_obuft_8_iopad (
            .OE(N__3740),
            .DIN(N__3739),
            .DOUT(N__3738),
            .PACKAGEPIN(p_vLED[8]));
    defparam p_vLED_obuft_8_preio.NEG_TRIGGER=1'b0;
    defparam p_vLED_obuft_8_preio.PIN_TYPE=6'b101001;
    PRE_IO p_vLED_obuft_8_preio (
            .PADOEN(N__3740),
            .PADOUT(N__3739),
            .PADIN(N__3738),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__2608),
            .DIN0(),
            .DOUT0(N__3071),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__830 (
            .O(N__3721),
            .I(N__3718));
    LocalMux I__829 (
            .O(N__3718),
            .I(p_hLED_cl_10_iZ0Z_0));
    IoInMux I__828 (
            .O(N__3715),
            .I(N__3712));
    LocalMux I__827 (
            .O(N__3712),
            .I(N__3709));
    Span4Mux_s1_h I__826 (
            .O(N__3709),
            .I(N__3706));
    Span4Mux_v I__825 (
            .O(N__3706),
            .I(N__3703));
    Odrv4 I__824 (
            .O(N__3703),
            .I(N_417_i));
    InMux I__823 (
            .O(N__3700),
            .I(N__3697));
    LocalMux I__822 (
            .O(N__3697),
            .I(N__3694));
    Odrv12 I__821 (
            .O(N__3694),
            .I(p_hLED_cl_9_iZ0Z_0));
    IoInMux I__820 (
            .O(N__3691),
            .I(N__3688));
    LocalMux I__819 (
            .O(N__3688),
            .I(N__3685));
    IoSpan4Mux I__818 (
            .O(N__3685),
            .I(N__3682));
    Span4Mux_s3_v I__817 (
            .O(N__3682),
            .I(N__3679));
    Odrv4 I__816 (
            .O(N__3679),
            .I(N_418_i));
    InMux I__815 (
            .O(N__3676),
            .I(N__3673));
    LocalMux I__814 (
            .O(N__3673),
            .I(N__3670));
    Span12Mux_s9_v I__813 (
            .O(N__3670),
            .I(N__3667));
    Odrv12 I__812 (
            .O(N__3667),
            .I(p_hLED_cl_1_iZ0Z_0));
    IoInMux I__811 (
            .O(N__3664),
            .I(N__3661));
    LocalMux I__810 (
            .O(N__3661),
            .I(N_413_i));
    InMux I__809 (
            .O(N__3658),
            .I(N__3655));
    LocalMux I__808 (
            .O(N__3655),
            .I(N__3652));
    Odrv12 I__807 (
            .O(N__3652),
            .I(p_hLED_cl_11_iZ0Z_0));
    IoInMux I__806 (
            .O(N__3649),
            .I(N__3646));
    LocalMux I__805 (
            .O(N__3646),
            .I(N__3643));
    Span4Mux_s0_h I__804 (
            .O(N__3643),
            .I(N__3640));
    Odrv4 I__803 (
            .O(N__3640),
            .I(N_420_i));
    InMux I__802 (
            .O(N__3637),
            .I(N__3634));
    LocalMux I__801 (
            .O(N__3634),
            .I(N__3631));
    Span4Mux_v I__800 (
            .O(N__3631),
            .I(N__3628));
    Odrv4 I__799 (
            .O(N__3628),
            .I(p_hLED_cl_12_iZ0Z_0));
    IoInMux I__798 (
            .O(N__3625),
            .I(N__3622));
    LocalMux I__797 (
            .O(N__3622),
            .I(N_415_i));
    InMux I__796 (
            .O(N__3619),
            .I(N__3616));
    LocalMux I__795 (
            .O(N__3616),
            .I(N__3613));
    Odrv12 I__794 (
            .O(N__3613),
            .I(p_hLED_cl_5_iZ0Z_0));
    IoInMux I__793 (
            .O(N__3610),
            .I(N__3607));
    LocalMux I__792 (
            .O(N__3607),
            .I(N_419_i));
    InMux I__791 (
            .O(N__3604),
            .I(N__3601));
    LocalMux I__790 (
            .O(N__3601),
            .I(p_hLED_cl_2_iZ0Z_0));
    IoInMux I__789 (
            .O(N__3598),
            .I(N__3595));
    LocalMux I__788 (
            .O(N__3595),
            .I(N_409_i));
    InMux I__787 (
            .O(N__3592),
            .I(N__3589));
    LocalMux I__786 (
            .O(N__3589),
            .I(p_hLED_cl_3_iZ0Z_0));
    CascadeMux I__785 (
            .O(N__3586),
            .I(N__3577));
    InMux I__784 (
            .O(N__3585),
            .I(N__3550));
    InMux I__783 (
            .O(N__3584),
            .I(N__3550));
    InMux I__782 (
            .O(N__3583),
            .I(N__3550));
    InMux I__781 (
            .O(N__3582),
            .I(N__3550));
    InMux I__780 (
            .O(N__3581),
            .I(N__3550));
    InMux I__779 (
            .O(N__3580),
            .I(N__3550));
    InMux I__778 (
            .O(N__3577),
            .I(N__3547));
    InMux I__777 (
            .O(N__3576),
            .I(N__3538));
    InMux I__776 (
            .O(N__3575),
            .I(N__3538));
    InMux I__775 (
            .O(N__3574),
            .I(N__3538));
    InMux I__774 (
            .O(N__3573),
            .I(N__3538));
    InMux I__773 (
            .O(N__3572),
            .I(N__3535));
    InMux I__772 (
            .O(N__3571),
            .I(N__3526));
    InMux I__771 (
            .O(N__3570),
            .I(N__3526));
    InMux I__770 (
            .O(N__3569),
            .I(N__3526));
    InMux I__769 (
            .O(N__3568),
            .I(N__3526));
    InMux I__768 (
            .O(N__3567),
            .I(N__3515));
    InMux I__767 (
            .O(N__3566),
            .I(N__3515));
    InMux I__766 (
            .O(N__3565),
            .I(N__3515));
    InMux I__765 (
            .O(N__3564),
            .I(N__3515));
    InMux I__764 (
            .O(N__3563),
            .I(N__3515));
    LocalMux I__763 (
            .O(N__3550),
            .I(N__3512));
    LocalMux I__762 (
            .O(N__3547),
            .I(N__3509));
    LocalMux I__761 (
            .O(N__3538),
            .I(N__3504));
    LocalMux I__760 (
            .O(N__3535),
            .I(N__3504));
    LocalMux I__759 (
            .O(N__3526),
            .I(hIndexZ0Z_3));
    LocalMux I__758 (
            .O(N__3515),
            .I(hIndexZ0Z_3));
    Odrv4 I__757 (
            .O(N__3512),
            .I(hIndexZ0Z_3));
    Odrv4 I__756 (
            .O(N__3509),
            .I(hIndexZ0Z_3));
    Odrv4 I__755 (
            .O(N__3504),
            .I(hIndexZ0Z_3));
    InMux I__754 (
            .O(N__3493),
            .I(N__3467));
    InMux I__753 (
            .O(N__3492),
            .I(N__3467));
    InMux I__752 (
            .O(N__3491),
            .I(N__3467));
    InMux I__751 (
            .O(N__3490),
            .I(N__3467));
    InMux I__750 (
            .O(N__3489),
            .I(N__3467));
    InMux I__749 (
            .O(N__3488),
            .I(N__3467));
    InMux I__748 (
            .O(N__3487),
            .I(N__3458));
    InMux I__747 (
            .O(N__3486),
            .I(N__3458));
    InMux I__746 (
            .O(N__3485),
            .I(N__3458));
    InMux I__745 (
            .O(N__3484),
            .I(N__3458));
    InMux I__744 (
            .O(N__3483),
            .I(N__3452));
    InMux I__743 (
            .O(N__3482),
            .I(N__3444));
    InMux I__742 (
            .O(N__3481),
            .I(N__3444));
    InMux I__741 (
            .O(N__3480),
            .I(N__3444));
    LocalMux I__740 (
            .O(N__3467),
            .I(N__3441));
    LocalMux I__739 (
            .O(N__3458),
            .I(N__3438));
    InMux I__738 (
            .O(N__3457),
            .I(N__3431));
    InMux I__737 (
            .O(N__3456),
            .I(N__3431));
    InMux I__736 (
            .O(N__3455),
            .I(N__3431));
    LocalMux I__735 (
            .O(N__3452),
            .I(N__3428));
    InMux I__734 (
            .O(N__3451),
            .I(N__3425));
    LocalMux I__733 (
            .O(N__3444),
            .I(hIndexZ0Z_2));
    Odrv4 I__732 (
            .O(N__3441),
            .I(hIndexZ0Z_2));
    Odrv4 I__731 (
            .O(N__3438),
            .I(hIndexZ0Z_2));
    LocalMux I__730 (
            .O(N__3431),
            .I(hIndexZ0Z_2));
    Odrv12 I__729 (
            .O(N__3428),
            .I(hIndexZ0Z_2));
    LocalMux I__728 (
            .O(N__3425),
            .I(hIndexZ0Z_2));
    CascadeMux I__727 (
            .O(N__3412),
            .I(N__3396));
    CascadeMux I__726 (
            .O(N__3411),
            .I(N__3393));
    CascadeMux I__725 (
            .O(N__3410),
            .I(N__3390));
    CascadeMux I__724 (
            .O(N__3409),
            .I(N__3387));
    CascadeMux I__723 (
            .O(N__3408),
            .I(N__3384));
    CascadeMux I__722 (
            .O(N__3407),
            .I(N__3381));
    CascadeMux I__721 (
            .O(N__3406),
            .I(N__3376));
    CascadeMux I__720 (
            .O(N__3405),
            .I(N__3373));
    CascadeMux I__719 (
            .O(N__3404),
            .I(N__3370));
    CascadeMux I__718 (
            .O(N__3403),
            .I(N__3367));
    CascadeMux I__717 (
            .O(N__3402),
            .I(N__3364));
    InMux I__716 (
            .O(N__3401),
            .I(N__3351));
    InMux I__715 (
            .O(N__3400),
            .I(N__3351));
    InMux I__714 (
            .O(N__3399),
            .I(N__3351));
    InMux I__713 (
            .O(N__3396),
            .I(N__3351));
    InMux I__712 (
            .O(N__3393),
            .I(N__3351));
    InMux I__711 (
            .O(N__3390),
            .I(N__3351));
    InMux I__710 (
            .O(N__3387),
            .I(N__3342));
    InMux I__709 (
            .O(N__3384),
            .I(N__3342));
    InMux I__708 (
            .O(N__3381),
            .I(N__3342));
    InMux I__707 (
            .O(N__3380),
            .I(N__3342));
    InMux I__706 (
            .O(N__3379),
            .I(N__3338));
    InMux I__705 (
            .O(N__3376),
            .I(N__3334));
    InMux I__704 (
            .O(N__3373),
            .I(N__3329));
    InMux I__703 (
            .O(N__3370),
            .I(N__3329));
    InMux I__702 (
            .O(N__3367),
            .I(N__3324));
    InMux I__701 (
            .O(N__3364),
            .I(N__3324));
    LocalMux I__700 (
            .O(N__3351),
            .I(N__3321));
    LocalMux I__699 (
            .O(N__3342),
            .I(N__3318));
    InMux I__698 (
            .O(N__3341),
            .I(N__3315));
    LocalMux I__697 (
            .O(N__3338),
            .I(N__3312));
    InMux I__696 (
            .O(N__3337),
            .I(N__3309));
    LocalMux I__695 (
            .O(N__3334),
            .I(hIndexZ0Z_1));
    LocalMux I__694 (
            .O(N__3329),
            .I(hIndexZ0Z_1));
    LocalMux I__693 (
            .O(N__3324),
            .I(hIndexZ0Z_1));
    Odrv4 I__692 (
            .O(N__3321),
            .I(hIndexZ0Z_1));
    Odrv4 I__691 (
            .O(N__3318),
            .I(hIndexZ0Z_1));
    LocalMux I__690 (
            .O(N__3315),
            .I(hIndexZ0Z_1));
    Odrv4 I__689 (
            .O(N__3312),
            .I(hIndexZ0Z_1));
    LocalMux I__688 (
            .O(N__3309),
            .I(hIndexZ0Z_1));
    CascadeMux I__687 (
            .O(N__3292),
            .I(N__3286));
    CascadeMux I__686 (
            .O(N__3291),
            .I(N__3277));
    CascadeMux I__685 (
            .O(N__3290),
            .I(N__3274));
    CascadeMux I__684 (
            .O(N__3289),
            .I(N__3271));
    InMux I__683 (
            .O(N__3286),
            .I(N__3262));
    InMux I__682 (
            .O(N__3285),
            .I(N__3262));
    InMux I__681 (
            .O(N__3284),
            .I(N__3262));
    InMux I__680 (
            .O(N__3283),
            .I(N__3262));
    InMux I__679 (
            .O(N__3282),
            .I(N__3249));
    InMux I__678 (
            .O(N__3281),
            .I(N__3249));
    InMux I__677 (
            .O(N__3280),
            .I(N__3249));
    InMux I__676 (
            .O(N__3277),
            .I(N__3249));
    InMux I__675 (
            .O(N__3274),
            .I(N__3249));
    InMux I__674 (
            .O(N__3271),
            .I(N__3249));
    LocalMux I__673 (
            .O(N__3262),
            .I(N__3234));
    LocalMux I__672 (
            .O(N__3249),
            .I(N__3234));
    InMux I__671 (
            .O(N__3248),
            .I(N__3231));
    InMux I__670 (
            .O(N__3247),
            .I(N__3225));
    InMux I__669 (
            .O(N__3246),
            .I(N__3225));
    InMux I__668 (
            .O(N__3245),
            .I(N__3220));
    InMux I__667 (
            .O(N__3244),
            .I(N__3220));
    InMux I__666 (
            .O(N__3243),
            .I(N__3213));
    InMux I__665 (
            .O(N__3242),
            .I(N__3213));
    InMux I__664 (
            .O(N__3241),
            .I(N__3213));
    InMux I__663 (
            .O(N__3240),
            .I(N__3210));
    InMux I__662 (
            .O(N__3239),
            .I(N__3207));
    Span4Mux_v I__661 (
            .O(N__3234),
            .I(N__3204));
    LocalMux I__660 (
            .O(N__3231),
            .I(N__3201));
    InMux I__659 (
            .O(N__3230),
            .I(N__3198));
    LocalMux I__658 (
            .O(N__3225),
            .I(hIndexZ0Z_0));
    LocalMux I__657 (
            .O(N__3220),
            .I(hIndexZ0Z_0));
    LocalMux I__656 (
            .O(N__3213),
            .I(hIndexZ0Z_0));
    LocalMux I__655 (
            .O(N__3210),
            .I(hIndexZ0Z_0));
    LocalMux I__654 (
            .O(N__3207),
            .I(hIndexZ0Z_0));
    Odrv4 I__653 (
            .O(N__3204),
            .I(hIndexZ0Z_0));
    Odrv4 I__652 (
            .O(N__3201),
            .I(hIndexZ0Z_0));
    LocalMux I__651 (
            .O(N__3198),
            .I(hIndexZ0Z_0));
    ClkMux I__650 (
            .O(N__3181),
            .I(N__3142));
    ClkMux I__649 (
            .O(N__3180),
            .I(N__3142));
    ClkMux I__648 (
            .O(N__3179),
            .I(N__3142));
    ClkMux I__647 (
            .O(N__3178),
            .I(N__3142));
    ClkMux I__646 (
            .O(N__3177),
            .I(N__3142));
    ClkMux I__645 (
            .O(N__3176),
            .I(N__3142));
    ClkMux I__644 (
            .O(N__3175),
            .I(N__3142));
    ClkMux I__643 (
            .O(N__3174),
            .I(N__3142));
    ClkMux I__642 (
            .O(N__3173),
            .I(N__3142));
    ClkMux I__641 (
            .O(N__3172),
            .I(N__3142));
    ClkMux I__640 (
            .O(N__3171),
            .I(N__3142));
    ClkMux I__639 (
            .O(N__3170),
            .I(N__3142));
    ClkMux I__638 (
            .O(N__3169),
            .I(N__3142));
    GlobalMux I__637 (
            .O(N__3142),
            .I(N__3139));
    gio2CtrlBuf I__636 (
            .O(N__3139),
            .I(p_clk12_c_g));
    CEMux I__635 (
            .O(N__3136),
            .I(N__3132));
    CEMux I__634 (
            .O(N__3135),
            .I(N__3128));
    LocalMux I__633 (
            .O(N__3132),
            .I(N__3125));
    CEMux I__632 (
            .O(N__3131),
            .I(N__3122));
    LocalMux I__631 (
            .O(N__3128),
            .I(N__3119));
    Span4Mux_v I__630 (
            .O(N__3125),
            .I(N__3114));
    LocalMux I__629 (
            .O(N__3122),
            .I(N__3114));
    Span4Mux_v I__628 (
            .O(N__3119),
            .I(N__3109));
    Span4Mux_s0_h I__627 (
            .O(N__3114),
            .I(N__3109));
    Span4Mux_h I__626 (
            .O(N__3109),
            .I(N__3106));
    Odrv4 I__625 (
            .O(N__3106),
            .I(p_hLED52));
    InMux I__624 (
            .O(N__3103),
            .I(N__3100));
    LocalMux I__623 (
            .O(N__3100),
            .I(p_hLED_cl_13_iZ0Z_0));
    IoInMux I__622 (
            .O(N__3097),
            .I(N__3094));
    LocalMux I__621 (
            .O(N__3094),
            .I(N__3091));
    Span4Mux_s0_h I__620 (
            .O(N__3091),
            .I(N__3088));
    Odrv4 I__619 (
            .O(N__3088),
            .I(N_416_i));
    InMux I__618 (
            .O(N__3085),
            .I(N__3082));
    LocalMux I__617 (
            .O(N__3082),
            .I(p_hLED_cl_8_iZ0Z_0));
    IoInMux I__616 (
            .O(N__3079),
            .I(N__3076));
    LocalMux I__615 (
            .O(N__3076),
            .I(N_411_i));
    IoInMux I__614 (
            .O(N__3073),
            .I(N__3067));
    IoInMux I__613 (
            .O(N__3072),
            .I(N__3064));
    IoInMux I__612 (
            .O(N__3071),
            .I(N__3059));
    IoInMux I__611 (
            .O(N__3070),
            .I(N__3056));
    LocalMux I__610 (
            .O(N__3067),
            .I(N__3051));
    LocalMux I__609 (
            .O(N__3064),
            .I(N__3051));
    IoInMux I__608 (
            .O(N__3063),
            .I(N__3048));
    IoInMux I__607 (
            .O(N__3062),
            .I(N__3045));
    LocalMux I__606 (
            .O(N__3059),
            .I(N__3038));
    LocalMux I__605 (
            .O(N__3056),
            .I(N__3038));
    IoSpan4Mux I__604 (
            .O(N__3051),
            .I(N__3038));
    LocalMux I__603 (
            .O(N__3048),
            .I(N__3035));
    LocalMux I__602 (
            .O(N__3045),
            .I(N__3032));
    Span4Mux_s0_h I__601 (
            .O(N__3038),
            .I(N__3025));
    Span4Mux_s0_h I__600 (
            .O(N__3035),
            .I(N__3020));
    Span4Mux_s0_h I__599 (
            .O(N__3032),
            .I(N__3020));
    IoInMux I__598 (
            .O(N__3031),
            .I(N__3017));
    IoInMux I__597 (
            .O(N__3030),
            .I(N__3014));
    IoInMux I__596 (
            .O(N__3029),
            .I(N__3011));
    IoInMux I__595 (
            .O(N__3028),
            .I(N__3008));
    Odrv4 I__594 (
            .O(N__3025),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__593 (
            .O(N__3020),
            .I(CONSTANT_ONE_NET));
    LocalMux I__592 (
            .O(N__3017),
            .I(CONSTANT_ONE_NET));
    LocalMux I__591 (
            .O(N__3014),
            .I(CONSTANT_ONE_NET));
    LocalMux I__590 (
            .O(N__3011),
            .I(CONSTANT_ONE_NET));
    LocalMux I__589 (
            .O(N__3008),
            .I(CONSTANT_ONE_NET));
    InMux I__588 (
            .O(N__2995),
            .I(N__2992));
    LocalMux I__587 (
            .O(N__2992),
            .I(N__2989));
    Span4Mux_v I__586 (
            .O(N__2989),
            .I(N__2986));
    Odrv4 I__585 (
            .O(N__2986),
            .I(p_hLED_cl_7_iZ0Z_0));
    InMux I__584 (
            .O(N__2983),
            .I(N__2980));
    LocalMux I__583 (
            .O(N__2980),
            .I(N__2977));
    Odrv4 I__582 (
            .O(N__2977),
            .I(p_hLED_cl_iZ0Z_0));
    InMux I__581 (
            .O(N__2974),
            .I(N__2967));
    InMux I__580 (
            .O(N__2973),
            .I(N__2967));
    InMux I__579 (
            .O(N__2972),
            .I(N__2964));
    LocalMux I__578 (
            .O(N__2967),
            .I(N_58));
    LocalMux I__577 (
            .O(N__2964),
            .I(N_58));
    InMux I__576 (
            .O(N__2959),
            .I(N__2956));
    LocalMux I__575 (
            .O(N__2956),
            .I(p_hLED_cl_14_iZ0Z_0));
    IoInMux I__574 (
            .O(N__2953),
            .I(N__2950));
    LocalMux I__573 (
            .O(N__2950),
            .I(N_406_i));
    InMux I__572 (
            .O(N__2947),
            .I(N__2944));
    LocalMux I__571 (
            .O(N__2944),
            .I(p_hLED_cl_4_iZ0Z_0));
    IoInMux I__570 (
            .O(N__2941),
            .I(N__2938));
    LocalMux I__569 (
            .O(N__2938),
            .I(N_408_i));
    IoInMux I__568 (
            .O(N__2935),
            .I(N__2932));
    LocalMux I__567 (
            .O(N__2932),
            .I(N_407_i));
    IoInMux I__566 (
            .O(N__2929),
            .I(N__2926));
    LocalMux I__565 (
            .O(N__2926),
            .I(N__2923));
    IoSpan4Mux I__564 (
            .O(N__2923),
            .I(N__2920));
    Span4Mux_s1_h I__563 (
            .O(N__2920),
            .I(N__2917));
    Odrv4 I__562 (
            .O(N__2917),
            .I(N_410_i));
    InMux I__561 (
            .O(N__2914),
            .I(N__2911));
    LocalMux I__560 (
            .O(N__2911),
            .I(p_hLED_cl_6_iZ0Z_0));
    InMux I__559 (
            .O(N__2908),
            .I(N__2905));
    LocalMux I__558 (
            .O(N__2905),
            .I(N__2902));
    Span4Mux_s3_v I__557 (
            .O(N__2902),
            .I(N__2899));
    Odrv4 I__556 (
            .O(N__2899),
            .I(p_vLED_cl_4_iZ0Z_0));
    IoInMux I__555 (
            .O(N__2896),
            .I(N__2893));
    LocalMux I__554 (
            .O(N__2893),
            .I(N_427_i));
    InMux I__553 (
            .O(N__2890),
            .I(N__2887));
    LocalMux I__552 (
            .O(N__2887),
            .I(N__2884));
    Span4Mux_s3_h I__551 (
            .O(N__2884),
            .I(N__2881));
    Odrv4 I__550 (
            .O(N__2881),
            .I(p_vLED_cl_7_iZ0Z_0));
    IoInMux I__549 (
            .O(N__2878),
            .I(N__2875));
    LocalMux I__548 (
            .O(N__2875),
            .I(N_426_i));
    IoInMux I__547 (
            .O(N__2872),
            .I(N__2869));
    LocalMux I__546 (
            .O(N__2869),
            .I(N__2866));
    Span4Mux_s3_v I__545 (
            .O(N__2866),
            .I(N__2863));
    Odrv4 I__544 (
            .O(N__2863),
            .I(N_414_i));
    InMux I__543 (
            .O(N__2860),
            .I(N__2857));
    LocalMux I__542 (
            .O(N__2857),
            .I(N__2854));
    Odrv12 I__541 (
            .O(N__2854),
            .I(p_vLED_cl_5_iZ0Z_0));
    IoInMux I__540 (
            .O(N__2851),
            .I(N__2848));
    LocalMux I__539 (
            .O(N__2848),
            .I(N__2845));
    Span4Mux_s0_h I__538 (
            .O(N__2845),
            .I(N__2842));
    Sp12to4 I__537 (
            .O(N__2842),
            .I(N__2839));
    Odrv12 I__536 (
            .O(N__2839),
            .I(N_421_i));
    CascadeMux I__535 (
            .O(N__2836),
            .I(N_58_cascade_));
    InMux I__534 (
            .O(N__2833),
            .I(N__2830));
    LocalMux I__533 (
            .O(N__2830),
            .I(N__2827));
    Span4Mux_v I__532 (
            .O(N__2827),
            .I(N__2824));
    Odrv4 I__531 (
            .O(N__2824),
            .I(p_vLED_cl_1_iZ0Z_0));
    IoInMux I__530 (
            .O(N__2821),
            .I(N__2818));
    LocalMux I__529 (
            .O(N__2818),
            .I(N__2815));
    Odrv12 I__528 (
            .O(N__2815),
            .I(N_423_i));
    InMux I__527 (
            .O(N__2812),
            .I(N__2807));
    InMux I__526 (
            .O(N__2811),
            .I(N__2804));
    InMux I__525 (
            .O(N__2810),
            .I(N__2801));
    LocalMux I__524 (
            .O(N__2807),
            .I(N__2798));
    LocalMux I__523 (
            .O(N__2804),
            .I(ballXZ0Z_1));
    LocalMux I__522 (
            .O(N__2801),
            .I(ballXZ0Z_1));
    Odrv12 I__521 (
            .O(N__2798),
            .I(ballXZ0Z_1));
    CascadeMux I__520 (
            .O(N__2791),
            .I(N__2787));
    CascadeMux I__519 (
            .O(N__2790),
            .I(N__2783));
    InMux I__518 (
            .O(N__2787),
            .I(N__2780));
    InMux I__517 (
            .O(N__2786),
            .I(N__2777));
    InMux I__516 (
            .O(N__2783),
            .I(N__2774));
    LocalMux I__515 (
            .O(N__2780),
            .I(N__2771));
    LocalMux I__514 (
            .O(N__2777),
            .I(ballXZ0Z_2));
    LocalMux I__513 (
            .O(N__2774),
            .I(ballXZ0Z_2));
    Odrv12 I__512 (
            .O(N__2771),
            .I(ballXZ0Z_2));
    InMux I__511 (
            .O(N__2764),
            .I(N__2759));
    InMux I__510 (
            .O(N__2763),
            .I(N__2754));
    InMux I__509 (
            .O(N__2762),
            .I(N__2754));
    LocalMux I__508 (
            .O(N__2759),
            .I(N__2751));
    LocalMux I__507 (
            .O(N__2754),
            .I(ballXZ0Z_0));
    Odrv12 I__506 (
            .O(N__2751),
            .I(ballXZ0Z_0));
    InMux I__505 (
            .O(N__2746),
            .I(N__2743));
    LocalMux I__504 (
            .O(N__2743),
            .I(p_hLED52_NE_0));
    InMux I__503 (
            .O(N__2740),
            .I(N__2737));
    LocalMux I__502 (
            .O(N__2737),
            .I(N_70_i));
    CascadeMux I__501 (
            .O(N__2734),
            .I(N__2731));
    InMux I__500 (
            .O(N__2731),
            .I(N__2728));
    LocalMux I__499 (
            .O(N__2728),
            .I(N__2723));
    InMux I__498 (
            .O(N__2727),
            .I(N__2718));
    InMux I__497 (
            .O(N__2726),
            .I(N__2718));
    Span4Mux_h I__496 (
            .O(N__2723),
            .I(N__2715));
    LocalMux I__495 (
            .O(N__2718),
            .I(ballXZ0Z_3));
    Odrv4 I__494 (
            .O(N__2715),
            .I(ballXZ0Z_3));
    InMux I__493 (
            .O(N__2710),
            .I(N__2706));
    InMux I__492 (
            .O(N__2709),
            .I(N__2703));
    LocalMux I__491 (
            .O(N__2706),
            .I(N__2700));
    LocalMux I__490 (
            .O(N__2703),
            .I(ctrZ0Z_15));
    Odrv4 I__489 (
            .O(N__2700),
            .I(ctrZ0Z_15));
    InMux I__488 (
            .O(N__2695),
            .I(ctr_cry_14));
    InMux I__487 (
            .O(N__2692),
            .I(N__2689));
    LocalMux I__486 (
            .O(N__2689),
            .I(N__2685));
    InMux I__485 (
            .O(N__2688),
            .I(N__2682));
    Span4Mux_h I__484 (
            .O(N__2685),
            .I(N__2679));
    LocalMux I__483 (
            .O(N__2682),
            .I(ctrZ0Z_16));
    Odrv4 I__482 (
            .O(N__2679),
            .I(ctrZ0Z_16));
    InMux I__481 (
            .O(N__2674),
            .I(bfn_9_9_0_));
    InMux I__480 (
            .O(N__2671),
            .I(N__2668));
    LocalMux I__479 (
            .O(N__2668),
            .I(N__2664));
    InMux I__478 (
            .O(N__2667),
            .I(N__2661));
    Span4Mux_h I__477 (
            .O(N__2664),
            .I(N__2658));
    LocalMux I__476 (
            .O(N__2661),
            .I(ctrZ0Z_17));
    Odrv4 I__475 (
            .O(N__2658),
            .I(ctrZ0Z_17));
    InMux I__474 (
            .O(N__2653),
            .I(ctr_cry_16));
    InMux I__473 (
            .O(N__2650),
            .I(ctr_cry_17));
    InMux I__472 (
            .O(N__2647),
            .I(N__2643));
    InMux I__471 (
            .O(N__2646),
            .I(N__2640));
    LocalMux I__470 (
            .O(N__2643),
            .I(N__2637));
    LocalMux I__469 (
            .O(N__2640),
            .I(ctrZ0Z_18));
    Odrv4 I__468 (
            .O(N__2637),
            .I(ctrZ0Z_18));
    IoInMux I__467 (
            .O(N__2632),
            .I(N__2629));
    LocalMux I__466 (
            .O(N__2629),
            .I(N__2626));
    Span4Mux_s1_v I__465 (
            .O(N__2626),
            .I(N__2623));
    Odrv4 I__464 (
            .O(N__2623),
            .I(N_412_i));
    InMux I__463 (
            .O(N__2620),
            .I(N__2617));
    LocalMux I__462 (
            .O(N__2617),
            .I(N__2614));
    Span4Mux_s3_v I__461 (
            .O(N__2614),
            .I(N__2611));
    Odrv4 I__460 (
            .O(N__2611),
            .I(p_vLED_cl_iZ0Z_0));
    IoInMux I__459 (
            .O(N__2608),
            .I(N__2605));
    LocalMux I__458 (
            .O(N__2605),
            .I(N__2602));
    Span4Mux_s1_h I__457 (
            .O(N__2602),
            .I(N__2599));
    Odrv4 I__456 (
            .O(N__2599),
            .I(N_429_i));
    InMux I__455 (
            .O(N__2596),
            .I(N__2593));
    LocalMux I__454 (
            .O(N__2593),
            .I(N__2590));
    Odrv4 I__453 (
            .O(N__2590),
            .I(p_vLED_cl_6_iZ0Z_0));
    IoInMux I__452 (
            .O(N__2587),
            .I(N__2584));
    LocalMux I__451 (
            .O(N__2584),
            .I(N__2581));
    Odrv4 I__450 (
            .O(N__2581),
            .I(N_425_i));
    InMux I__449 (
            .O(N__2578),
            .I(N__2575));
    LocalMux I__448 (
            .O(N__2575),
            .I(N__2572));
    Odrv4 I__447 (
            .O(N__2572),
            .I(p_vLED_cl_8_iZ0Z_0));
    IoInMux I__446 (
            .O(N__2569),
            .I(N__2566));
    LocalMux I__445 (
            .O(N__2566),
            .I(N__2563));
    Odrv12 I__444 (
            .O(N__2563),
            .I(N_424_i));
    InMux I__443 (
            .O(N__2560),
            .I(N__2557));
    LocalMux I__442 (
            .O(N__2557),
            .I(N__2554));
    Odrv4 I__441 (
            .O(N__2554),
            .I(p_vLED_cl_3_iZ0Z_0));
    IoInMux I__440 (
            .O(N__2551),
            .I(N__2548));
    LocalMux I__439 (
            .O(N__2548),
            .I(N__2545));
    IoSpan4Mux I__438 (
            .O(N__2545),
            .I(N__2542));
    Odrv4 I__437 (
            .O(N__2542),
            .I(N_422_i));
    CascadeMux I__436 (
            .O(N__2539),
            .I(N__2535));
    InMux I__435 (
            .O(N__2538),
            .I(N__2532));
    InMux I__434 (
            .O(N__2535),
            .I(N__2529));
    LocalMux I__433 (
            .O(N__2532),
            .I(N__2524));
    LocalMux I__432 (
            .O(N__2529),
            .I(N__2524));
    Odrv4 I__431 (
            .O(N__2524),
            .I(ctrZ0Z_7));
    InMux I__430 (
            .O(N__2521),
            .I(ctr_cry_6));
    InMux I__429 (
            .O(N__2518),
            .I(N__2514));
    InMux I__428 (
            .O(N__2517),
            .I(N__2511));
    LocalMux I__427 (
            .O(N__2514),
            .I(ctrZ0Z_8));
    LocalMux I__426 (
            .O(N__2511),
            .I(ctrZ0Z_8));
    InMux I__425 (
            .O(N__2506),
            .I(bfn_9_8_0_));
    InMux I__424 (
            .O(N__2503),
            .I(N__2499));
    InMux I__423 (
            .O(N__2502),
            .I(N__2496));
    LocalMux I__422 (
            .O(N__2499),
            .I(N__2493));
    LocalMux I__421 (
            .O(N__2496),
            .I(ctrZ0Z_9));
    Odrv4 I__420 (
            .O(N__2493),
            .I(ctrZ0Z_9));
    InMux I__419 (
            .O(N__2488),
            .I(ctr_cry_8));
    InMux I__418 (
            .O(N__2485),
            .I(N__2481));
    InMux I__417 (
            .O(N__2484),
            .I(N__2478));
    LocalMux I__416 (
            .O(N__2481),
            .I(ctrZ0Z_10));
    LocalMux I__415 (
            .O(N__2478),
            .I(ctrZ0Z_10));
    InMux I__414 (
            .O(N__2473),
            .I(ctr_cry_9));
    InMux I__413 (
            .O(N__2470),
            .I(N__2466));
    InMux I__412 (
            .O(N__2469),
            .I(N__2463));
    LocalMux I__411 (
            .O(N__2466),
            .I(ctrZ0Z_11));
    LocalMux I__410 (
            .O(N__2463),
            .I(ctrZ0Z_11));
    InMux I__409 (
            .O(N__2458),
            .I(ctr_cry_10));
    InMux I__408 (
            .O(N__2455),
            .I(N__2451));
    InMux I__407 (
            .O(N__2454),
            .I(N__2448));
    LocalMux I__406 (
            .O(N__2451),
            .I(ctrZ0Z_12));
    LocalMux I__405 (
            .O(N__2448),
            .I(ctrZ0Z_12));
    InMux I__404 (
            .O(N__2443),
            .I(ctr_cry_11));
    InMux I__403 (
            .O(N__2440),
            .I(N__2436));
    InMux I__402 (
            .O(N__2439),
            .I(N__2433));
    LocalMux I__401 (
            .O(N__2436),
            .I(ctrZ0Z_13));
    LocalMux I__400 (
            .O(N__2433),
            .I(ctrZ0Z_13));
    InMux I__399 (
            .O(N__2428),
            .I(ctr_cry_12));
    CascadeMux I__398 (
            .O(N__2425),
            .I(N__2421));
    InMux I__397 (
            .O(N__2424),
            .I(N__2418));
    InMux I__396 (
            .O(N__2421),
            .I(N__2415));
    LocalMux I__395 (
            .O(N__2418),
            .I(ctrZ0Z_14));
    LocalMux I__394 (
            .O(N__2415),
            .I(ctrZ0Z_14));
    InMux I__393 (
            .O(N__2410),
            .I(ctr_cry_13));
    InMux I__392 (
            .O(N__2407),
            .I(N__2401));
    InMux I__391 (
            .O(N__2406),
            .I(N__2398));
    InMux I__390 (
            .O(N__2405),
            .I(N__2395));
    InMux I__389 (
            .O(N__2404),
            .I(N__2392));
    LocalMux I__388 (
            .O(N__2401),
            .I(p_vLED33));
    LocalMux I__387 (
            .O(N__2398),
            .I(p_vLED33));
    LocalMux I__386 (
            .O(N__2395),
            .I(p_vLED33));
    LocalMux I__385 (
            .O(N__2392),
            .I(p_vLED33));
    CascadeMux I__384 (
            .O(N__2383),
            .I(N_57_i_cascade_));
    CascadeMux I__383 (
            .O(N__2380),
            .I(N__2377));
    InMux I__382 (
            .O(N__2377),
            .I(N__2373));
    InMux I__381 (
            .O(N__2376),
            .I(N__2370));
    LocalMux I__380 (
            .O(N__2373),
            .I(N_76));
    LocalMux I__379 (
            .O(N__2370),
            .I(N_76));
    InMux I__378 (
            .O(N__2365),
            .I(N__2346));
    InMux I__377 (
            .O(N__2364),
            .I(N__2346));
    InMux I__376 (
            .O(N__2363),
            .I(N__2346));
    InMux I__375 (
            .O(N__2362),
            .I(N__2346));
    InMux I__374 (
            .O(N__2361),
            .I(N__2346));
    InMux I__373 (
            .O(N__2360),
            .I(N__2346));
    CascadeMux I__372 (
            .O(N__2359),
            .I(N__2340));
    LocalMux I__371 (
            .O(N__2346),
            .I(N__2335));
    InMux I__370 (
            .O(N__2345),
            .I(N__2328));
    InMux I__369 (
            .O(N__2344),
            .I(N__2328));
    InMux I__368 (
            .O(N__2343),
            .I(N__2328));
    InMux I__367 (
            .O(N__2340),
            .I(N__2325));
    InMux I__366 (
            .O(N__2339),
            .I(N__2320));
    InMux I__365 (
            .O(N__2338),
            .I(N__2320));
    Odrv4 I__364 (
            .O(N__2335),
            .I(vIndexZ0Z_0));
    LocalMux I__363 (
            .O(N__2328),
            .I(vIndexZ0Z_0));
    LocalMux I__362 (
            .O(N__2325),
            .I(vIndexZ0Z_0));
    LocalMux I__361 (
            .O(N__2320),
            .I(vIndexZ0Z_0));
    InMux I__360 (
            .O(N__2311),
            .I(N__2307));
    InMux I__359 (
            .O(N__2310),
            .I(N__2304));
    LocalMux I__358 (
            .O(N__2307),
            .I(N__2299));
    LocalMux I__357 (
            .O(N__2304),
            .I(N__2299));
    Odrv4 I__356 (
            .O(N__2299),
            .I(ctrZ0Z_0));
    InMux I__355 (
            .O(N__2296),
            .I(bfn_9_7_0_));
    CascadeMux I__354 (
            .O(N__2293),
            .I(N__2289));
    InMux I__353 (
            .O(N__2292),
            .I(N__2286));
    InMux I__352 (
            .O(N__2289),
            .I(N__2283));
    LocalMux I__351 (
            .O(N__2286),
            .I(ctrZ0Z_1));
    LocalMux I__350 (
            .O(N__2283),
            .I(ctrZ0Z_1));
    InMux I__349 (
            .O(N__2278),
            .I(ctr_cry_0));
    InMux I__348 (
            .O(N__2275),
            .I(N__2271));
    InMux I__347 (
            .O(N__2274),
            .I(N__2268));
    LocalMux I__346 (
            .O(N__2271),
            .I(ctrZ0Z_2));
    LocalMux I__345 (
            .O(N__2268),
            .I(ctrZ0Z_2));
    InMux I__344 (
            .O(N__2263),
            .I(ctr_cry_1));
    InMux I__343 (
            .O(N__2260),
            .I(N__2256));
    InMux I__342 (
            .O(N__2259),
            .I(N__2253));
    LocalMux I__341 (
            .O(N__2256),
            .I(ctrZ0Z_3));
    LocalMux I__340 (
            .O(N__2253),
            .I(ctrZ0Z_3));
    InMux I__339 (
            .O(N__2248),
            .I(ctr_cry_2));
    InMux I__338 (
            .O(N__2245),
            .I(N__2241));
    InMux I__337 (
            .O(N__2244),
            .I(N__2238));
    LocalMux I__336 (
            .O(N__2241),
            .I(ctrZ0Z_4));
    LocalMux I__335 (
            .O(N__2238),
            .I(ctrZ0Z_4));
    InMux I__334 (
            .O(N__2233),
            .I(ctr_cry_3));
    InMux I__333 (
            .O(N__2230),
            .I(N__2226));
    InMux I__332 (
            .O(N__2229),
            .I(N__2223));
    LocalMux I__331 (
            .O(N__2226),
            .I(ctrZ0Z_5));
    LocalMux I__330 (
            .O(N__2223),
            .I(ctrZ0Z_5));
    InMux I__329 (
            .O(N__2218),
            .I(ctr_cry_4));
    CascadeMux I__328 (
            .O(N__2215),
            .I(N__2211));
    InMux I__327 (
            .O(N__2214),
            .I(N__2208));
    InMux I__326 (
            .O(N__2211),
            .I(N__2205));
    LocalMux I__325 (
            .O(N__2208),
            .I(ctrZ0Z_6));
    LocalMux I__324 (
            .O(N__2205),
            .I(ctrZ0Z_6));
    InMux I__323 (
            .O(N__2200),
            .I(ctr_cry_5));
    InMux I__322 (
            .O(N__2197),
            .I(N__2194));
    LocalMux I__321 (
            .O(N__2194),
            .I(N__2191));
    Odrv4 I__320 (
            .O(N__2191),
            .I(p_vLED_cl_2_iZ0Z_0));
    InMux I__319 (
            .O(N__2188),
            .I(N__2185));
    LocalMux I__318 (
            .O(N__2185),
            .I(N__2182));
    Odrv12 I__317 (
            .O(N__2182),
            .I(p_vLED_cl_9_iZ0Z_0));
    CEMux I__316 (
            .O(N__2179),
            .I(N__2175));
    CEMux I__315 (
            .O(N__2178),
            .I(N__2172));
    LocalMux I__314 (
            .O(N__2175),
            .I(N__2169));
    LocalMux I__313 (
            .O(N__2172),
            .I(N__2166));
    Odrv4 I__312 (
            .O(N__2169),
            .I(p_vLED37));
    Odrv4 I__311 (
            .O(N__2166),
            .I(p_vLED37));
    InMux I__310 (
            .O(N__2161),
            .I(N__2141));
    InMux I__309 (
            .O(N__2160),
            .I(N__2141));
    InMux I__308 (
            .O(N__2159),
            .I(N__2141));
    InMux I__307 (
            .O(N__2158),
            .I(N__2141));
    InMux I__306 (
            .O(N__2157),
            .I(N__2141));
    InMux I__305 (
            .O(N__2156),
            .I(N__2141));
    CascadeMux I__304 (
            .O(N__2155),
            .I(N__2135));
    InMux I__303 (
            .O(N__2154),
            .I(N__2131));
    LocalMux I__302 (
            .O(N__2141),
            .I(N__2128));
    InMux I__301 (
            .O(N__2140),
            .I(N__2121));
    InMux I__300 (
            .O(N__2139),
            .I(N__2121));
    InMux I__299 (
            .O(N__2138),
            .I(N__2121));
    InMux I__298 (
            .O(N__2135),
            .I(N__2116));
    InMux I__297 (
            .O(N__2134),
            .I(N__2116));
    LocalMux I__296 (
            .O(N__2131),
            .I(N__2113));
    Odrv4 I__295 (
            .O(N__2128),
            .I(vIndexZ0Z_2));
    LocalMux I__294 (
            .O(N__2121),
            .I(vIndexZ0Z_2));
    LocalMux I__293 (
            .O(N__2116),
            .I(vIndexZ0Z_2));
    Odrv4 I__292 (
            .O(N__2113),
            .I(vIndexZ0Z_2));
    CascadeMux I__291 (
            .O(N__2104),
            .I(N__2097));
    CascadeMux I__290 (
            .O(N__2103),
            .I(N__2094));
    CascadeMux I__289 (
            .O(N__2102),
            .I(N__2091));
    CascadeMux I__288 (
            .O(N__2101),
            .I(N__2085));
    CascadeMux I__287 (
            .O(N__2100),
            .I(N__2082));
    InMux I__286 (
            .O(N__2097),
            .I(N__2068));
    InMux I__285 (
            .O(N__2094),
            .I(N__2068));
    InMux I__284 (
            .O(N__2091),
            .I(N__2068));
    InMux I__283 (
            .O(N__2090),
            .I(N__2068));
    InMux I__282 (
            .O(N__2089),
            .I(N__2068));
    InMux I__281 (
            .O(N__2088),
            .I(N__2068));
    InMux I__280 (
            .O(N__2085),
            .I(N__2058));
    InMux I__279 (
            .O(N__2082),
            .I(N__2058));
    InMux I__278 (
            .O(N__2081),
            .I(N__2058));
    LocalMux I__277 (
            .O(N__2068),
            .I(N__2055));
    InMux I__276 (
            .O(N__2067),
            .I(N__2052));
    InMux I__275 (
            .O(N__2066),
            .I(N__2049));
    InMux I__274 (
            .O(N__2065),
            .I(N__2046));
    LocalMux I__273 (
            .O(N__2058),
            .I(vIndexZ0Z_1));
    Odrv4 I__272 (
            .O(N__2055),
            .I(vIndexZ0Z_1));
    LocalMux I__271 (
            .O(N__2052),
            .I(vIndexZ0Z_1));
    LocalMux I__270 (
            .O(N__2049),
            .I(vIndexZ0Z_1));
    LocalMux I__269 (
            .O(N__2046),
            .I(vIndexZ0Z_1));
    CascadeMux I__268 (
            .O(N__2035),
            .I(N__2027));
    CascadeMux I__267 (
            .O(N__2034),
            .I(N__2024));
    CascadeMux I__266 (
            .O(N__2033),
            .I(N__2021));
    InMux I__265 (
            .O(N__2032),
            .I(N__2006));
    InMux I__264 (
            .O(N__2031),
            .I(N__2006));
    InMux I__263 (
            .O(N__2030),
            .I(N__2006));
    InMux I__262 (
            .O(N__2027),
            .I(N__2006));
    InMux I__261 (
            .O(N__2024),
            .I(N__2006));
    InMux I__260 (
            .O(N__2021),
            .I(N__2006));
    CascadeMux I__259 (
            .O(N__2020),
            .I(N__2001));
    CascadeMux I__258 (
            .O(N__2019),
            .I(N__1996));
    LocalMux I__257 (
            .O(N__2006),
            .I(N__1993));
    InMux I__256 (
            .O(N__2005),
            .I(N__1986));
    InMux I__255 (
            .O(N__2004),
            .I(N__1986));
    InMux I__254 (
            .O(N__2001),
            .I(N__1986));
    InMux I__253 (
            .O(N__2000),
            .I(N__1983));
    InMux I__252 (
            .O(N__1999),
            .I(N__1980));
    InMux I__251 (
            .O(N__1996),
            .I(N__1977));
    Odrv4 I__250 (
            .O(N__1993),
            .I(vIndexZ0Z_3));
    LocalMux I__249 (
            .O(N__1986),
            .I(vIndexZ0Z_3));
    LocalMux I__248 (
            .O(N__1983),
            .I(vIndexZ0Z_3));
    LocalMux I__247 (
            .O(N__1980),
            .I(vIndexZ0Z_3));
    LocalMux I__246 (
            .O(N__1977),
            .I(vIndexZ0Z_3));
    CascadeMux I__245 (
            .O(N__1966),
            .I(N_76_cascade_));
    InMux I__244 (
            .O(N__1963),
            .I(N__1960));
    LocalMux I__243 (
            .O(N__1960),
            .I(N_57_i));
    CascadeMux I__242 (
            .O(N__1957),
            .I(ballXVel12_10_cascade_));
    InMux I__241 (
            .O(N__1954),
            .I(N__1951));
    LocalMux I__240 (
            .O(N__1951),
            .I(ballXVel12_12));
    CascadeMux I__239 (
            .O(N__1948),
            .I(ballXVel12_14_cascade_));
    InMux I__238 (
            .O(N__1945),
            .I(N__1942));
    LocalMux I__237 (
            .O(N__1942),
            .I(ballXVel12_11));
    CascadeMux I__236 (
            .O(N__1939),
            .I(N__1933));
    CascadeMux I__235 (
            .O(N__1938),
            .I(N__1928));
    CascadeMux I__234 (
            .O(N__1937),
            .I(N__1922));
    InMux I__233 (
            .O(N__1936),
            .I(N__1918));
    InMux I__232 (
            .O(N__1933),
            .I(N__1913));
    InMux I__231 (
            .O(N__1932),
            .I(N__1913));
    InMux I__230 (
            .O(N__1931),
            .I(N__1904));
    InMux I__229 (
            .O(N__1928),
            .I(N__1904));
    InMux I__228 (
            .O(N__1927),
            .I(N__1904));
    InMux I__227 (
            .O(N__1926),
            .I(N__1904));
    InMux I__226 (
            .O(N__1925),
            .I(N__1897));
    InMux I__225 (
            .O(N__1922),
            .I(N__1897));
    InMux I__224 (
            .O(N__1921),
            .I(N__1897));
    LocalMux I__223 (
            .O(N__1918),
            .I(ballXVel12));
    LocalMux I__222 (
            .O(N__1913),
            .I(ballXVel12));
    LocalMux I__221 (
            .O(N__1904),
            .I(ballXVel12));
    LocalMux I__220 (
            .O(N__1897),
            .I(ballXVel12));
    InMux I__219 (
            .O(N__1888),
            .I(N__1885));
    LocalMux I__218 (
            .O(N__1885),
            .I(ballXVel12_13));
    IoInMux I__217 (
            .O(N__1882),
            .I(N__1879));
    LocalMux I__216 (
            .O(N__1879),
            .I(N__1876));
    Odrv12 I__215 (
            .O(N__1876),
            .I(N_430_i));
    IoInMux I__214 (
            .O(N__1873),
            .I(N__1870));
    LocalMux I__213 (
            .O(N__1870),
            .I(N__1867));
    Odrv12 I__212 (
            .O(N__1867),
            .I(N_428_i));
    InMux I__211 (
            .O(N__1864),
            .I(N__1861));
    LocalMux I__210 (
            .O(N__1861),
            .I(N_67_i));
    InMux I__209 (
            .O(N__1858),
            .I(un1_vIndex_2_cry_0));
    InMux I__208 (
            .O(N__1855),
            .I(un1_vIndex_2_cry_1));
    InMux I__207 (
            .O(N__1852),
            .I(un1_vIndex_2_cry_2));
    InMux I__206 (
            .O(N__1849),
            .I(N__1844));
    InMux I__205 (
            .O(N__1848),
            .I(N__1839));
    InMux I__204 (
            .O(N__1847),
            .I(N__1839));
    LocalMux I__203 (
            .O(N__1844),
            .I(ballYZ0Z_0));
    LocalMux I__202 (
            .O(N__1839),
            .I(ballYZ0Z_0));
    CascadeMux I__201 (
            .O(N__1834),
            .I(N__1831));
    InMux I__200 (
            .O(N__1831),
            .I(N__1826));
    InMux I__199 (
            .O(N__1830),
            .I(N__1823));
    InMux I__198 (
            .O(N__1829),
            .I(N__1820));
    LocalMux I__197 (
            .O(N__1826),
            .I(ballYZ0Z_1));
    LocalMux I__196 (
            .O(N__1823),
            .I(ballYZ0Z_1));
    LocalMux I__195 (
            .O(N__1820),
            .I(ballYZ0Z_1));
    CascadeMux I__194 (
            .O(N__1813),
            .I(ballYVel_s_1_0_0_cascade_));
    InMux I__193 (
            .O(N__1810),
            .I(N__1803));
    InMux I__192 (
            .O(N__1809),
            .I(N__1798));
    InMux I__191 (
            .O(N__1808),
            .I(N__1798));
    InMux I__190 (
            .O(N__1807),
            .I(N__1793));
    InMux I__189 (
            .O(N__1806),
            .I(N__1793));
    LocalMux I__188 (
            .O(N__1803),
            .I(ballYVelZ0Z_0));
    LocalMux I__187 (
            .O(N__1798),
            .I(ballYVelZ0Z_0));
    LocalMux I__186 (
            .O(N__1793),
            .I(ballYVelZ0Z_0));
    CascadeMux I__185 (
            .O(N__1786),
            .I(N__1782));
    InMux I__184 (
            .O(N__1785),
            .I(N__1778));
    InMux I__183 (
            .O(N__1782),
            .I(N__1773));
    InMux I__182 (
            .O(N__1781),
            .I(N__1773));
    LocalMux I__181 (
            .O(N__1778),
            .I(ballYZ0Z_2));
    LocalMux I__180 (
            .O(N__1773),
            .I(ballYZ0Z_2));
    CascadeMux I__179 (
            .O(N__1768),
            .I(N__1764));
    CascadeMux I__178 (
            .O(N__1767),
            .I(N__1760));
    InMux I__177 (
            .O(N__1764),
            .I(N__1757));
    InMux I__176 (
            .O(N__1763),
            .I(N__1752));
    InMux I__175 (
            .O(N__1760),
            .I(N__1752));
    LocalMux I__174 (
            .O(N__1757),
            .I(N__1747));
    LocalMux I__173 (
            .O(N__1752),
            .I(N__1747));
    Odrv4 I__172 (
            .O(N__1747),
            .I(ballYZ0Z_3));
    InMux I__171 (
            .O(N__1744),
            .I(N__1741));
    LocalMux I__170 (
            .O(N__1741),
            .I(p_vLED37_NE_0));
    InMux I__169 (
            .O(N__1738),
            .I(un1_ballX_3_cry_0));
    InMux I__168 (
            .O(N__1735),
            .I(un1_ballX_3_cry_1));
    InMux I__167 (
            .O(N__1732),
            .I(un1_ballX_3_cry_2));
    CascadeMux I__166 (
            .O(N__1729),
            .I(ballXVel_s_1_0_0_cascade_));
    CascadeMux I__165 (
            .O(N__1726),
            .I(N__1723));
    InMux I__164 (
            .O(N__1723),
            .I(N__1720));
    LocalMux I__163 (
            .O(N__1720),
            .I(ballXVel_RNIFI1J4_0Z0Z_0));
    InMux I__162 (
            .O(N__1717),
            .I(N__1702));
    InMux I__161 (
            .O(N__1716),
            .I(N__1702));
    InMux I__160 (
            .O(N__1715),
            .I(N__1702));
    InMux I__159 (
            .O(N__1714),
            .I(N__1702));
    InMux I__158 (
            .O(N__1713),
            .I(N__1702));
    LocalMux I__157 (
            .O(N__1702),
            .I(ballXVelZ0Z_0));
    CascadeMux I__156 (
            .O(N__1699),
            .I(N__1696));
    InMux I__155 (
            .O(N__1696),
            .I(N__1693));
    LocalMux I__154 (
            .O(N__1693),
            .I(ballXVel_RNIFI1J4Z0Z_0));
    InMux I__153 (
            .O(N__1690),
            .I(un1_ballY_4_cry_0));
    InMux I__152 (
            .O(N__1687),
            .I(un1_ballY_4_cry_1));
    InMux I__151 (
            .O(N__1684),
            .I(un1_ballY_4_cry_2));
    CascadeMux I__150 (
            .O(N__1681),
            .I(N__1678));
    InMux I__149 (
            .O(N__1678),
            .I(N__1675));
    LocalMux I__148 (
            .O(N__1675),
            .I(ballYVel_RNIGOGN4_0Z0Z_0));
    CascadeMux I__147 (
            .O(N__1672),
            .I(N__1669));
    InMux I__146 (
            .O(N__1669),
            .I(N__1666));
    LocalMux I__145 (
            .O(N__1666),
            .I(ballYVel_RNIGOGN4Z0Z_0));
    defparam IN_MUX_bfv_9_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_7_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(ctr_cry_7),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(ctr_cry_15),
            .carryinitout(bfn_9_9_0_));
    defparam IN_MUX_bfv_7_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_6_0_));
    defparam IN_MUX_bfv_8_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_6_0_));
    defparam IN_MUX_bfv_7_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_7_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam ballY_0_LC_7_6_0.C_ON=1'b1;
    defparam ballY_0_LC_7_6_0.SEQ_MODE=4'b1000;
    defparam ballY_0_LC_7_6_0.LUT_INIT=16'b0011110000111100;
    LogicCell40 ballY_0_LC_7_6_0 (
            .in0(_gnd_net_),
            .in1(N__1849),
            .in2(N__1938),
            .in3(_gnd_net_),
            .lcout(ballYZ0Z_0),
            .ltout(),
            .carryin(bfn_7_6_0_),
            .carryout(un1_ballY_4_cry_0),
            .clk(N__3171),
            .ce(),
            .sr(_gnd_net_));
    defparam ballY_1_LC_7_6_1.C_ON=1'b1;
    defparam ballY_1_LC_7_6_1.SEQ_MODE=4'b1000;
    defparam ballY_1_LC_7_6_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 ballY_1_LC_7_6_1 (
            .in0(_gnd_net_),
            .in1(N__1830),
            .in2(N__1672),
            .in3(N__1690),
            .lcout(ballYZ0Z_1),
            .ltout(),
            .carryin(un1_ballY_4_cry_0),
            .carryout(un1_ballY_4_cry_1),
            .clk(N__3171),
            .ce(),
            .sr(_gnd_net_));
    defparam ballY_2_LC_7_6_2.C_ON=1'b1;
    defparam ballY_2_LC_7_6_2.SEQ_MODE=4'b1000;
    defparam ballY_2_LC_7_6_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 ballY_2_LC_7_6_2 (
            .in0(_gnd_net_),
            .in1(N__1785),
            .in2(N__1681),
            .in3(N__1687),
            .lcout(ballYZ0Z_2),
            .ltout(),
            .carryin(un1_ballY_4_cry_1),
            .carryout(un1_ballY_4_cry_2),
            .clk(N__3171),
            .ce(),
            .sr(_gnd_net_));
    defparam ballY_3_LC_7_6_3.C_ON=1'b0;
    defparam ballY_3_LC_7_6_3.SEQ_MODE=4'b1000;
    defparam ballY_3_LC_7_6_3.LUT_INIT=16'b1000011101111000;
    LogicCell40 ballY_3_LC_7_6_3 (
            .in0(N__1810),
            .in1(N__1931),
            .in2(N__1768),
            .in3(N__1684),
            .lcout(ballYZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3171),
            .ce(),
            .sr(_gnd_net_));
    defparam ballYVel_RNIGOGN4_0_0_LC_7_6_5.C_ON=1'b0;
    defparam ballYVel_RNIGOGN4_0_0_LC_7_6_5.SEQ_MODE=4'b0000;
    defparam ballYVel_RNIGOGN4_0_0_LC_7_6_5.LUT_INIT=16'b1100110000000000;
    LogicCell40 ballYVel_RNIGOGN4_0_0_LC_7_6_5 (
            .in0(_gnd_net_),
            .in1(N__1807),
            .in2(_gnd_net_),
            .in3(N__1927),
            .lcout(ballYVel_RNIGOGN4_0Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ballYVel_RNIGOGN4_0_LC_7_6_7.C_ON=1'b0;
    defparam ballYVel_RNIGOGN4_0_LC_7_6_7.SEQ_MODE=4'b0000;
    defparam ballYVel_RNIGOGN4_0_LC_7_6_7.LUT_INIT=16'b1100110000000000;
    LogicCell40 ballYVel_RNIGOGN4_0_LC_7_6_7 (
            .in0(_gnd_net_),
            .in1(N__1806),
            .in2(_gnd_net_),
            .in3(N__1926),
            .lcout(ballYVel_RNIGOGN4Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ballX_0_LC_7_7_0.C_ON=1'b1;
    defparam ballX_0_LC_7_7_0.SEQ_MODE=4'b1000;
    defparam ballX_0_LC_7_7_0.LUT_INIT=16'b0011110000111100;
    LogicCell40 ballX_0_LC_7_7_0 (
            .in0(_gnd_net_),
            .in1(N__2762),
            .in2(N__1937),
            .in3(_gnd_net_),
            .lcout(ballXZ0Z_0),
            .ltout(),
            .carryin(bfn_7_7_0_),
            .carryout(un1_ballX_3_cry_0),
            .clk(N__3169),
            .ce(),
            .sr(_gnd_net_));
    defparam ballX_1_LC_7_7_1.C_ON=1'b1;
    defparam ballX_1_LC_7_7_1.SEQ_MODE=4'b1000;
    defparam ballX_1_LC_7_7_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 ballX_1_LC_7_7_1 (
            .in0(_gnd_net_),
            .in1(N__2811),
            .in2(N__1699),
            .in3(N__1738),
            .lcout(ballXZ0Z_1),
            .ltout(),
            .carryin(un1_ballX_3_cry_0),
            .carryout(un1_ballX_3_cry_1),
            .clk(N__3169),
            .ce(),
            .sr(_gnd_net_));
    defparam ballX_2_LC_7_7_2.C_ON=1'b1;
    defparam ballX_2_LC_7_7_2.SEQ_MODE=4'b1000;
    defparam ballX_2_LC_7_7_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 ballX_2_LC_7_7_2 (
            .in0(_gnd_net_),
            .in1(N__2786),
            .in2(N__1726),
            .in3(N__1735),
            .lcout(ballXZ0Z_2),
            .ltout(),
            .carryin(un1_ballX_3_cry_1),
            .carryout(un1_ballX_3_cry_2),
            .clk(N__3169),
            .ce(),
            .sr(_gnd_net_));
    defparam ballX_3_LC_7_7_3.C_ON=1'b0;
    defparam ballX_3_LC_7_7_3.SEQ_MODE=4'b1000;
    defparam ballX_3_LC_7_7_3.LUT_INIT=16'b1001010101101010;
    LogicCell40 ballX_3_LC_7_7_3 (
            .in0(N__2726),
            .in1(N__1717),
            .in2(N__1939),
            .in3(N__1732),
            .lcout(ballXZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3169),
            .ce(),
            .sr(_gnd_net_));
    defparam ballXVel_RNO_0_0_LC_7_7_4.C_ON=1'b0;
    defparam ballXVel_RNO_0_0_LC_7_7_4.SEQ_MODE=4'b0000;
    defparam ballXVel_RNO_0_0_LC_7_7_4.LUT_INIT=16'b0001001000000000;
    LogicCell40 ballXVel_RNO_0_0_LC_7_7_4 (
            .in0(N__1715),
            .in1(N__2810),
            .in2(N__2790),
            .in3(N__2763),
            .lcout(),
            .ltout(ballXVel_s_1_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ballXVel_0_LC_7_7_5.C_ON=1'b0;
    defparam ballXVel_0_LC_7_7_5.SEQ_MODE=4'b1000;
    defparam ballXVel_0_LC_7_7_5.LUT_INIT=16'b1010110011001100;
    LogicCell40 ballXVel_0_LC_7_7_5 (
            .in0(N__2727),
            .in1(N__1716),
            .in2(N__1729),
            .in3(N__1925),
            .lcout(ballXVelZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3169),
            .ce(),
            .sr(_gnd_net_));
    defparam ballXVel_RNIFI1J4_0_0_LC_7_7_6.C_ON=1'b0;
    defparam ballXVel_RNIFI1J4_0_0_LC_7_7_6.SEQ_MODE=4'b0000;
    defparam ballXVel_RNIFI1J4_0_0_LC_7_7_6.LUT_INIT=16'b1010101000000000;
    LogicCell40 ballXVel_RNIFI1J4_0_0_LC_7_7_6 (
            .in0(N__1714),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1932),
            .lcout(ballXVel_RNIFI1J4_0Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ballXVel_RNIFI1J4_0_LC_7_7_7.C_ON=1'b0;
    defparam ballXVel_RNIFI1J4_0_LC_7_7_7.SEQ_MODE=4'b0000;
    defparam ballXVel_RNIFI1J4_0_LC_7_7_7.LUT_INIT=16'b1100110000000000;
    LogicCell40 ballXVel_RNIFI1J4_0_LC_7_7_7 (
            .in0(_gnd_net_),
            .in1(N__1713),
            .in2(_gnd_net_),
            .in3(N__1921),
            .lcout(ballXVel_RNIFI1J4Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ballY_RNIKQR82_1_LC_8_5_3.C_ON=1'b0;
    defparam ballY_RNIKQR82_1_LC_8_5_3.SEQ_MODE=4'b0000;
    defparam ballY_RNIKQR82_1_LC_8_5_3.LUT_INIT=16'b0010000000000010;
    LogicCell40 ballY_RNIKQR82_1_LC_8_5_3 (
            .in0(N__1744),
            .in1(N__1864),
            .in2(N__1834),
            .in3(N__2066),
            .lcout(p_vLED37),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ballY_RNIIR6I_0_LC_8_6_0.C_ON=1'b1;
    defparam ballY_RNIIR6I_0_LC_8_6_0.SEQ_MODE=4'b0000;
    defparam ballY_RNIIR6I_0_LC_8_6_0.LUT_INIT=16'b0000111111110000;
    LogicCell40 ballY_RNIIR6I_0_LC_8_6_0 (
            .in0(_gnd_net_),
            .in1(N__1963),
            .in2(N__2359),
            .in3(N__1847),
            .lcout(N_67_i),
            .ltout(),
            .carryin(bfn_8_6_0_),
            .carryout(un1_vIndex_2_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam vIndex_1_LC_8_6_1.C_ON=1'b1;
    defparam vIndex_1_LC_8_6_1.SEQ_MODE=4'b1000;
    defparam vIndex_1_LC_8_6_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 vIndex_1_LC_8_6_1 (
            .in0(_gnd_net_),
            .in1(N__2067),
            .in2(_gnd_net_),
            .in3(N__1858),
            .lcout(vIndexZ0Z_1),
            .ltout(),
            .carryin(un1_vIndex_2_cry_0),
            .carryout(un1_vIndex_2_cry_1),
            .clk(N__3172),
            .ce(),
            .sr(_gnd_net_));
    defparam vIndex_2_LC_8_6_2.C_ON=1'b1;
    defparam vIndex_2_LC_8_6_2.SEQ_MODE=4'b1000;
    defparam vIndex_2_LC_8_6_2.LUT_INIT=16'b1010010101011010;
    LogicCell40 vIndex_2_LC_8_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2155),
            .in3(N__1855),
            .lcout(vIndexZ0Z_2),
            .ltout(),
            .carryin(un1_vIndex_2_cry_1),
            .carryout(un1_vIndex_2_cry_2),
            .clk(N__3172),
            .ce(),
            .sr(_gnd_net_));
    defparam vIndex_3_LC_8_6_3.C_ON=1'b0;
    defparam vIndex_3_LC_8_6_3.SEQ_MODE=4'b1000;
    defparam vIndex_3_LC_8_6_3.LUT_INIT=16'b0101000110100010;
    LogicCell40 vIndex_3_LC_8_6_3 (
            .in0(N__2000),
            .in1(N__2406),
            .in2(N__2380),
            .in3(N__1852),
            .lcout(vIndexZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3172),
            .ce(),
            .sr(_gnd_net_));
    defparam ballYVel_RNO_0_0_LC_8_6_5.C_ON=1'b0;
    defparam ballYVel_RNO_0_0_LC_8_6_5.SEQ_MODE=4'b0000;
    defparam ballYVel_RNO_0_0_LC_8_6_5.LUT_INIT=16'b0000001000000001;
    LogicCell40 ballYVel_RNO_0_0_LC_8_6_5 (
            .in0(N__1848),
            .in1(N__1829),
            .in2(N__1786),
            .in3(N__1808),
            .lcout(),
            .ltout(ballYVel_s_1_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ballYVel_0_LC_8_6_6.C_ON=1'b0;
    defparam ballYVel_0_LC_8_6_6.SEQ_MODE=4'b1000;
    defparam ballYVel_0_LC_8_6_6.LUT_INIT=16'b1100101010101010;
    LogicCell40 ballYVel_0_LC_8_6_6 (
            .in0(N__1809),
            .in1(N__1763),
            .in2(N__1813),
            .in3(N__1936),
            .lcout(ballYVelZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3172),
            .ce(),
            .sr(_gnd_net_));
    defparam ballY_RNIE1E41_3_LC_8_6_7.C_ON=1'b0;
    defparam ballY_RNIE1E41_3_LC_8_6_7.SEQ_MODE=4'b0000;
    defparam ballY_RNIE1E41_3_LC_8_6_7.LUT_INIT=16'b1000001001000001;
    LogicCell40 ballY_RNIE1E41_3_LC_8_6_7 (
            .in0(N__1781),
            .in1(N__1999),
            .in2(N__1767),
            .in3(N__2134),
            .lcout(p_vLED37_NE_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_RNIDIAM_7_LC_8_7_0.C_ON=1'b0;
    defparam ctr_RNIDIAM_7_LC_8_7_0.SEQ_MODE=4'b0000;
    defparam ctr_RNIDIAM_7_LC_8_7_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 ctr_RNIDIAM_7_LC_8_7_0 (
            .in0(N__2503),
            .in1(N__2517),
            .in2(N__2539),
            .in3(N__2484),
            .lcout(ballXVel12_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_RNIM4UE_3_LC_8_7_2.C_ON=1'b0;
    defparam ctr_RNIM4UE_3_LC_8_7_2.SEQ_MODE=4'b0000;
    defparam ctr_RNIM4UE_3_LC_8_7_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 ctr_RNIM4UE_3_LC_8_7_2 (
            .in0(N__2229),
            .in1(N__2244),
            .in2(N__2215),
            .in3(N__2259),
            .lcout(ballXVel12_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_RNI05AM_18_LC_8_7_3.C_ON=1'b0;
    defparam ctr_RNI05AM_18_LC_8_7_3.SEQ_MODE=4'b0000;
    defparam ctr_RNI05AM_18_LC_8_7_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 ctr_RNI05AM_18_LC_8_7_3 (
            .in0(N__2310),
            .in1(N__2647),
            .in2(N__2293),
            .in3(N__2274),
            .lcout(),
            .ltout(ballXVel12_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_RNIOJLN1_15_LC_8_7_4.C_ON=1'b0;
    defparam ctr_RNIOJLN1_15_LC_8_7_4.SEQ_MODE=4'b0000;
    defparam ctr_RNIOJLN1_15_LC_8_7_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 ctr_RNIOJLN1_15_LC_8_7_4 (
            .in0(N__2671),
            .in1(N__2692),
            .in2(N__1957),
            .in3(N__2710),
            .lcout(),
            .ltout(ballXVel12_14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_RNID5D94_3_LC_8_7_5.C_ON=1'b0;
    defparam ctr_RNID5D94_3_LC_8_7_5.SEQ_MODE=4'b0000;
    defparam ctr_RNID5D94_3_LC_8_7_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 ctr_RNID5D94_3_LC_8_7_5 (
            .in0(N__1888),
            .in1(N__1954),
            .in2(N__1948),
            .in3(N__1945),
            .lcout(ballXVel12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_RNIIQEC1_11_LC_8_8_0.C_ON=1'b0;
    defparam ctr_RNIIQEC1_11_LC_8_8_0.SEQ_MODE=4'b0000;
    defparam ctr_RNIIQEC1_11_LC_8_8_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 ctr_RNIIQEC1_11_LC_8_8_0 (
            .in0(N__2439),
            .in1(N__2454),
            .in2(N__2425),
            .in3(N__2469),
            .lcout(ballXVel12_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam p_vLED_obuft_RNO_9_LC_9_1_2.C_ON=1'b0;
    defparam p_vLED_obuft_RNO_9_LC_9_1_2.SEQ_MODE=4'b0000;
    defparam p_vLED_obuft_RNO_9_LC_9_1_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 p_vLED_obuft_RNO_9_LC_9_1_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2188),
            .lcout(N_430_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam p_vLED_obuft_RNO_7_LC_9_2_4.C_ON=1'b0;
    defparam p_vLED_obuft_RNO_7_LC_9_2_4.SEQ_MODE=4'b0000;
    defparam p_vLED_obuft_RNO_7_LC_9_2_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 p_vLED_obuft_RNO_7_LC_9_2_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2197),
            .lcout(N_428_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam p_vLED_cl_4_i_0_LC_9_4_1.C_ON=1'b0;
    defparam p_vLED_cl_4_i_0_LC_9_4_1.SEQ_MODE=4'b1000;
    defparam p_vLED_cl_4_i_0_LC_9_4_1.LUT_INIT=16'b1111111111110111;
    LogicCell40 p_vLED_cl_4_i_0_LC_9_4_1 (
            .in0(N__2157),
            .in1(N__2089),
            .in2(N__2034),
            .in3(N__2361),
            .lcout(p_vLED_cl_4_iZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3181),
            .ce(N__2179),
            .sr(_gnd_net_));
    defparam p_vLED_cl_i_0_LC_9_4_2.C_ON=1'b0;
    defparam p_vLED_cl_i_0_LC_9_4_2.SEQ_MODE=4'b1000;
    defparam p_vLED_cl_i_0_LC_9_4_2.LUT_INIT=16'b1111111111111011;
    LogicCell40 p_vLED_cl_i_0_LC_9_4_2 (
            .in0(N__2365),
            .in1(N__2032),
            .in2(N__2104),
            .in3(N__2161),
            .lcout(p_vLED_cl_iZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3181),
            .ce(N__2179),
            .sr(_gnd_net_));
    defparam p_vLED_cl_7_i_0_LC_9_4_4.C_ON=1'b0;
    defparam p_vLED_cl_7_i_0_LC_9_4_4.SEQ_MODE=4'b1000;
    defparam p_vLED_cl_7_i_0_LC_9_4_4.LUT_INIT=16'b1111110111111111;
    LogicCell40 p_vLED_cl_7_i_0_LC_9_4_4 (
            .in0(N__2363),
            .in1(N__2030),
            .in2(N__2102),
            .in3(N__2159),
            .lcout(p_vLED_cl_7_iZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3181),
            .ce(N__2179),
            .sr(_gnd_net_));
    defparam p_vLED_cl_2_i_0_LC_9_4_5.C_ON=1'b0;
    defparam p_vLED_cl_2_i_0_LC_9_4_5.SEQ_MODE=4'b1000;
    defparam p_vLED_cl_2_i_0_LC_9_4_5.LUT_INIT=16'b1111011111111111;
    LogicCell40 p_vLED_cl_2_i_0_LC_9_4_5 (
            .in0(N__2156),
            .in1(N__2088),
            .in2(N__2033),
            .in3(N__2360),
            .lcout(p_vLED_cl_2_iZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3181),
            .ce(N__2179),
            .sr(_gnd_net_));
    defparam p_vLED_cl_8_i_0_LC_9_4_6.C_ON=1'b0;
    defparam p_vLED_cl_8_i_0_LC_9_4_6.SEQ_MODE=4'b1000;
    defparam p_vLED_cl_8_i_0_LC_9_4_6.LUT_INIT=16'b1111111111011111;
    LogicCell40 p_vLED_cl_8_i_0_LC_9_4_6 (
            .in0(N__2364),
            .in1(N__2031),
            .in2(N__2103),
            .in3(N__2160),
            .lcout(p_vLED_cl_8_iZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3181),
            .ce(N__2179),
            .sr(_gnd_net_));
    defparam p_vLED_cl_6_i_0_LC_9_4_7.C_ON=1'b0;
    defparam p_vLED_cl_6_i_0_LC_9_4_7.SEQ_MODE=4'b1000;
    defparam p_vLED_cl_6_i_0_LC_9_4_7.LUT_INIT=16'b1111111111111101;
    LogicCell40 p_vLED_cl_6_i_0_LC_9_4_7 (
            .in0(N__2158),
            .in1(N__2090),
            .in2(N__2035),
            .in3(N__2362),
            .lcout(p_vLED_cl_6_iZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3181),
            .ce(N__2179),
            .sr(_gnd_net_));
    defparam p_vLED_cl_1_i_0_LC_9_5_1.C_ON=1'b0;
    defparam p_vLED_cl_1_i_0_LC_9_5_1.SEQ_MODE=4'b1000;
    defparam p_vLED_cl_1_i_0_LC_9_5_1.LUT_INIT=16'b1111111111111011;
    LogicCell40 p_vLED_cl_1_i_0_LC_9_5_1 (
            .in0(N__2138),
            .in1(N__2081),
            .in2(N__2020),
            .in3(N__2343),
            .lcout(p_vLED_cl_1_iZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3177),
            .ce(N__2178),
            .sr(_gnd_net_));
    defparam p_vLED_cl_9_i_0_LC_9_5_3.C_ON=1'b0;
    defparam p_vLED_cl_9_i_0_LC_9_5_3.SEQ_MODE=4'b1000;
    defparam p_vLED_cl_9_i_0_LC_9_5_3.LUT_INIT=16'b0011001100110011;
    LogicCell40 p_vLED_cl_9_i_0_LC_9_5_3 (
            .in0(_gnd_net_),
            .in1(N__2405),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(p_vLED_cl_9_iZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3177),
            .ce(N__2178),
            .sr(_gnd_net_));
    defparam p_vLED_cl_5_i_0_LC_9_5_4.C_ON=1'b0;
    defparam p_vLED_cl_5_i_0_LC_9_5_4.SEQ_MODE=4'b1000;
    defparam p_vLED_cl_5_i_0_LC_9_5_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 p_vLED_cl_5_i_0_LC_9_5_4 (
            .in0(N__2345),
            .in1(N__2140),
            .in2(N__2101),
            .in3(N__2005),
            .lcout(p_vLED_cl_5_iZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3177),
            .ce(N__2178),
            .sr(_gnd_net_));
    defparam p_vLED_cl_3_i_0_LC_9_5_6.C_ON=1'b0;
    defparam p_vLED_cl_3_i_0_LC_9_5_6.SEQ_MODE=4'b1000;
    defparam p_vLED_cl_3_i_0_LC_9_5_6.LUT_INIT=16'b1111111111111101;
    LogicCell40 p_vLED_cl_3_i_0_LC_9_5_6 (
            .in0(N__2344),
            .in1(N__2139),
            .in2(N__2100),
            .in3(N__2004),
            .lcout(p_vLED_cl_3_iZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3177),
            .ce(N__2178),
            .sr(_gnd_net_));
    defparam vIndex_RNIUK6M_3_LC_9_6_0.C_ON=1'b0;
    defparam vIndex_RNIUK6M_3_LC_9_6_0.SEQ_MODE=4'b0000;
    defparam vIndex_RNIUK6M_3_LC_9_6_0.LUT_INIT=16'b0001000000000000;
    LogicCell40 vIndex_RNIUK6M_3_LC_9_6_0 (
            .in0(N__2154),
            .in1(N__2065),
            .in2(N__2019),
            .in3(N__2338),
            .lcout(p_vLED33),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam hIndex_RNI6JO41_1_LC_9_6_1.C_ON=1'b0;
    defparam hIndex_RNI6JO41_1_LC_9_6_1.SEQ_MODE=4'b0000;
    defparam hIndex_RNI6JO41_1_LC_9_6_1.LUT_INIT=16'b1101111111111111;
    LogicCell40 hIndex_RNI6JO41_1_LC_9_6_1 (
            .in0(N__3483),
            .in1(N__3248),
            .in2(N__3586),
            .in3(N__3379),
            .lcout(N_76),
            .ltout(N_76_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam vIndex_RNI48VQ1_3_LC_9_6_2.C_ON=1'b0;
    defparam vIndex_RNI48VQ1_3_LC_9_6_2.SEQ_MODE=4'b0000;
    defparam vIndex_RNI48VQ1_3_LC_9_6_2.LUT_INIT=16'b0000000000001111;
    LogicCell40 vIndex_RNI48VQ1_3_LC_9_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1966),
            .in3(N__2404),
            .lcout(N_57_i),
            .ltout(N_57_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam vIndex_0_LC_9_6_3.C_ON=1'b0;
    defparam vIndex_0_LC_9_6_3.SEQ_MODE=4'b1000;
    defparam vIndex_0_LC_9_6_3.LUT_INIT=16'b0101101000010010;
    LogicCell40 vIndex_0_LC_9_6_3 (
            .in0(N__2339),
            .in1(N__2407),
            .in2(N__2383),
            .in3(N__2376),
            .lcout(vIndexZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3175),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_0_LC_9_7_0.C_ON=1'b1;
    defparam ctr_0_LC_9_7_0.SEQ_MODE=4'b1000;
    defparam ctr_0_LC_9_7_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_0_LC_9_7_0 (
            .in0(_gnd_net_),
            .in1(N__2311),
            .in2(_gnd_net_),
            .in3(N__2296),
            .lcout(ctrZ0Z_0),
            .ltout(),
            .carryin(bfn_9_7_0_),
            .carryout(ctr_cry_0),
            .clk(N__3173),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_1_LC_9_7_1.C_ON=1'b1;
    defparam ctr_1_LC_9_7_1.SEQ_MODE=4'b1000;
    defparam ctr_1_LC_9_7_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_1_LC_9_7_1 (
            .in0(_gnd_net_),
            .in1(N__2292),
            .in2(_gnd_net_),
            .in3(N__2278),
            .lcout(ctrZ0Z_1),
            .ltout(),
            .carryin(ctr_cry_0),
            .carryout(ctr_cry_1),
            .clk(N__3173),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_2_LC_9_7_2.C_ON=1'b1;
    defparam ctr_2_LC_9_7_2.SEQ_MODE=4'b1000;
    defparam ctr_2_LC_9_7_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_2_LC_9_7_2 (
            .in0(_gnd_net_),
            .in1(N__2275),
            .in2(_gnd_net_),
            .in3(N__2263),
            .lcout(ctrZ0Z_2),
            .ltout(),
            .carryin(ctr_cry_1),
            .carryout(ctr_cry_2),
            .clk(N__3173),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_3_LC_9_7_3.C_ON=1'b1;
    defparam ctr_3_LC_9_7_3.SEQ_MODE=4'b1000;
    defparam ctr_3_LC_9_7_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_3_LC_9_7_3 (
            .in0(_gnd_net_),
            .in1(N__2260),
            .in2(_gnd_net_),
            .in3(N__2248),
            .lcout(ctrZ0Z_3),
            .ltout(),
            .carryin(ctr_cry_2),
            .carryout(ctr_cry_3),
            .clk(N__3173),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_4_LC_9_7_4.C_ON=1'b1;
    defparam ctr_4_LC_9_7_4.SEQ_MODE=4'b1000;
    defparam ctr_4_LC_9_7_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_4_LC_9_7_4 (
            .in0(_gnd_net_),
            .in1(N__2245),
            .in2(_gnd_net_),
            .in3(N__2233),
            .lcout(ctrZ0Z_4),
            .ltout(),
            .carryin(ctr_cry_3),
            .carryout(ctr_cry_4),
            .clk(N__3173),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_5_LC_9_7_5.C_ON=1'b1;
    defparam ctr_5_LC_9_7_5.SEQ_MODE=4'b1000;
    defparam ctr_5_LC_9_7_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_5_LC_9_7_5 (
            .in0(_gnd_net_),
            .in1(N__2230),
            .in2(_gnd_net_),
            .in3(N__2218),
            .lcout(ctrZ0Z_5),
            .ltout(),
            .carryin(ctr_cry_4),
            .carryout(ctr_cry_5),
            .clk(N__3173),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_6_LC_9_7_6.C_ON=1'b1;
    defparam ctr_6_LC_9_7_6.SEQ_MODE=4'b1000;
    defparam ctr_6_LC_9_7_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_6_LC_9_7_6 (
            .in0(_gnd_net_),
            .in1(N__2214),
            .in2(_gnd_net_),
            .in3(N__2200),
            .lcout(ctrZ0Z_6),
            .ltout(),
            .carryin(ctr_cry_5),
            .carryout(ctr_cry_6),
            .clk(N__3173),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_7_LC_9_7_7.C_ON=1'b1;
    defparam ctr_7_LC_9_7_7.SEQ_MODE=4'b1000;
    defparam ctr_7_LC_9_7_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_7_LC_9_7_7 (
            .in0(_gnd_net_),
            .in1(N__2538),
            .in2(_gnd_net_),
            .in3(N__2521),
            .lcout(ctrZ0Z_7),
            .ltout(),
            .carryin(ctr_cry_6),
            .carryout(ctr_cry_7),
            .clk(N__3173),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_8_LC_9_8_0.C_ON=1'b1;
    defparam ctr_8_LC_9_8_0.SEQ_MODE=4'b1000;
    defparam ctr_8_LC_9_8_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_8_LC_9_8_0 (
            .in0(_gnd_net_),
            .in1(N__2518),
            .in2(_gnd_net_),
            .in3(N__2506),
            .lcout(ctrZ0Z_8),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(ctr_cry_8),
            .clk(N__3170),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_9_LC_9_8_1.C_ON=1'b1;
    defparam ctr_9_LC_9_8_1.SEQ_MODE=4'b1000;
    defparam ctr_9_LC_9_8_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_9_LC_9_8_1 (
            .in0(_gnd_net_),
            .in1(N__2502),
            .in2(_gnd_net_),
            .in3(N__2488),
            .lcout(ctrZ0Z_9),
            .ltout(),
            .carryin(ctr_cry_8),
            .carryout(ctr_cry_9),
            .clk(N__3170),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_10_LC_9_8_2.C_ON=1'b1;
    defparam ctr_10_LC_9_8_2.SEQ_MODE=4'b1000;
    defparam ctr_10_LC_9_8_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_10_LC_9_8_2 (
            .in0(_gnd_net_),
            .in1(N__2485),
            .in2(_gnd_net_),
            .in3(N__2473),
            .lcout(ctrZ0Z_10),
            .ltout(),
            .carryin(ctr_cry_9),
            .carryout(ctr_cry_10),
            .clk(N__3170),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_11_LC_9_8_3.C_ON=1'b1;
    defparam ctr_11_LC_9_8_3.SEQ_MODE=4'b1000;
    defparam ctr_11_LC_9_8_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_11_LC_9_8_3 (
            .in0(_gnd_net_),
            .in1(N__2470),
            .in2(_gnd_net_),
            .in3(N__2458),
            .lcout(ctrZ0Z_11),
            .ltout(),
            .carryin(ctr_cry_10),
            .carryout(ctr_cry_11),
            .clk(N__3170),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_12_LC_9_8_4.C_ON=1'b1;
    defparam ctr_12_LC_9_8_4.SEQ_MODE=4'b1000;
    defparam ctr_12_LC_9_8_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_12_LC_9_8_4 (
            .in0(_gnd_net_),
            .in1(N__2455),
            .in2(_gnd_net_),
            .in3(N__2443),
            .lcout(ctrZ0Z_12),
            .ltout(),
            .carryin(ctr_cry_11),
            .carryout(ctr_cry_12),
            .clk(N__3170),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_13_LC_9_8_5.C_ON=1'b1;
    defparam ctr_13_LC_9_8_5.SEQ_MODE=4'b1000;
    defparam ctr_13_LC_9_8_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_13_LC_9_8_5 (
            .in0(_gnd_net_),
            .in1(N__2440),
            .in2(_gnd_net_),
            .in3(N__2428),
            .lcout(ctrZ0Z_13),
            .ltout(),
            .carryin(ctr_cry_12),
            .carryout(ctr_cry_13),
            .clk(N__3170),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_14_LC_9_8_6.C_ON=1'b1;
    defparam ctr_14_LC_9_8_6.SEQ_MODE=4'b1000;
    defparam ctr_14_LC_9_8_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_14_LC_9_8_6 (
            .in0(_gnd_net_),
            .in1(N__2424),
            .in2(_gnd_net_),
            .in3(N__2410),
            .lcout(ctrZ0Z_14),
            .ltout(),
            .carryin(ctr_cry_13),
            .carryout(ctr_cry_14),
            .clk(N__3170),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_15_LC_9_8_7.C_ON=1'b1;
    defparam ctr_15_LC_9_8_7.SEQ_MODE=4'b1000;
    defparam ctr_15_LC_9_8_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_15_LC_9_8_7 (
            .in0(_gnd_net_),
            .in1(N__2709),
            .in2(_gnd_net_),
            .in3(N__2695),
            .lcout(ctrZ0Z_15),
            .ltout(),
            .carryin(ctr_cry_14),
            .carryout(ctr_cry_15),
            .clk(N__3170),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_16_LC_9_9_0.C_ON=1'b1;
    defparam ctr_16_LC_9_9_0.SEQ_MODE=4'b1000;
    defparam ctr_16_LC_9_9_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_16_LC_9_9_0 (
            .in0(_gnd_net_),
            .in1(N__2688),
            .in2(_gnd_net_),
            .in3(N__2674),
            .lcout(ctrZ0Z_16),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(ctr_cry_16),
            .clk(N__3174),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_17_LC_9_9_1.C_ON=1'b1;
    defparam ctr_17_LC_9_9_1.SEQ_MODE=4'b1000;
    defparam ctr_17_LC_9_9_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_17_LC_9_9_1 (
            .in0(_gnd_net_),
            .in1(N__2667),
            .in2(_gnd_net_),
            .in3(N__2653),
            .lcout(ctrZ0Z_17),
            .ltout(),
            .carryin(ctr_cry_16),
            .carryout(ctr_cry_17),
            .clk(N__3174),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_18_LC_9_9_2.C_ON=1'b0;
    defparam ctr_18_LC_9_9_2.SEQ_MODE=4'b1000;
    defparam ctr_18_LC_9_9_2.LUT_INIT=16'b0011001111001100;
    LogicCell40 ctr_18_LC_9_9_2 (
            .in0(_gnd_net_),
            .in1(N__2646),
            .in2(_gnd_net_),
            .in3(N__2650),
            .lcout(ctrZ0Z_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3174),
            .ce(),
            .sr(_gnd_net_));
    defparam p_hLED_obuft_RNO_6_LC_11_2_1.C_ON=1'b0;
    defparam p_hLED_obuft_RNO_6_LC_11_2_1.SEQ_MODE=4'b0000;
    defparam p_hLED_obuft_RNO_6_LC_11_2_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 p_hLED_obuft_RNO_6_LC_11_2_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2995),
            .lcout(N_412_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam p_vLED_obuft_RNO_8_LC_11_2_7.C_ON=1'b0;
    defparam p_vLED_obuft_RNO_8_LC_11_2_7.SEQ_MODE=4'b0000;
    defparam p_vLED_obuft_RNO_8_LC_11_2_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 p_vLED_obuft_RNO_8_LC_11_2_7 (
            .in0(N__2620),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_429_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam p_vLED_obuft_RNO_4_LC_11_4_3.C_ON=1'b0;
    defparam p_vLED_obuft_RNO_4_LC_11_4_3.SEQ_MODE=4'b0000;
    defparam p_vLED_obuft_RNO_4_LC_11_4_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 p_vLED_obuft_RNO_4_LC_11_4_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2596),
            .lcout(N_425_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam p_vLED_obuft_RNO_3_LC_11_4_5.C_ON=1'b0;
    defparam p_vLED_obuft_RNO_3_LC_11_4_5.SEQ_MODE=4'b0000;
    defparam p_vLED_obuft_RNO_3_LC_11_4_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 p_vLED_obuft_RNO_3_LC_11_4_5 (
            .in0(N__2578),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_424_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam p_vLED_obuft_RNO_1_LC_11_5_0.C_ON=1'b0;
    defparam p_vLED_obuft_RNO_1_LC_11_5_0.SEQ_MODE=4'b0000;
    defparam p_vLED_obuft_RNO_1_LC_11_5_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 p_vLED_obuft_RNO_1_LC_11_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2560),
            .lcout(N_422_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam hIndex_RNIJ9CI_1_LC_11_6_0.C_ON=1'b0;
    defparam hIndex_RNIJ9CI_1_LC_11_6_0.SEQ_MODE=4'b0000;
    defparam hIndex_RNIJ9CI_1_LC_11_6_0.LUT_INIT=16'b0011001111111111;
    LogicCell40 hIndex_RNIJ9CI_1_LC_11_6_0 (
            .in0(_gnd_net_),
            .in1(N__3341),
            .in2(_gnd_net_),
            .in3(N__3455),
            .lcout(N_58),
            .ltout(N_58_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam hIndex_0_LC_11_6_1.C_ON=1'b0;
    defparam hIndex_0_LC_11_6_1.SEQ_MODE=4'b1000;
    defparam hIndex_0_LC_11_6_1.LUT_INIT=16'b0011000000110011;
    LogicCell40 hIndex_0_LC_11_6_1 (
            .in0(_gnd_net_),
            .in1(N__3239),
            .in2(N__2836),
            .in3(N__3570),
            .lcout(hIndexZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3178),
            .ce(),
            .sr(_gnd_net_));
    defparam hIndex_1_LC_11_6_2.C_ON=1'b0;
    defparam hIndex_1_LC_11_6_2.SEQ_MODE=4'b1000;
    defparam hIndex_1_LC_11_6_2.LUT_INIT=16'b0000111101110000;
    LogicCell40 hIndex_1_LC_11_6_2 (
            .in0(N__3568),
            .in1(N__3456),
            .in2(N__3402),
            .in3(N__3244),
            .lcout(hIndexZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3178),
            .ce(),
            .sr(_gnd_net_));
    defparam hIndex_3_LC_11_6_3.C_ON=1'b0;
    defparam hIndex_3_LC_11_6_3.SEQ_MODE=4'b1000;
    defparam hIndex_3_LC_11_6_3.LUT_INIT=16'b1100110000100010;
    LogicCell40 hIndex_3_LC_11_6_3 (
            .in0(N__3240),
            .in1(N__2972),
            .in2(_gnd_net_),
            .in3(N__3571),
            .lcout(hIndexZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3178),
            .ce(),
            .sr(_gnd_net_));
    defparam hIndex_2_LC_11_6_4.C_ON=1'b0;
    defparam hIndex_2_LC_11_6_4.SEQ_MODE=4'b1000;
    defparam hIndex_2_LC_11_6_4.LUT_INIT=16'b0011110001001100;
    LogicCell40 hIndex_2_LC_11_6_4 (
            .in0(N__3569),
            .in1(N__3457),
            .in2(N__3403),
            .in3(N__3245),
            .lcout(hIndexZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3178),
            .ce(),
            .sr(_gnd_net_));
    defparam p_vLED_obuft_RNO_2_LC_11_6_5.C_ON=1'b0;
    defparam p_vLED_obuft_RNO_2_LC_11_6_5.SEQ_MODE=4'b0000;
    defparam p_vLED_obuft_RNO_2_LC_11_6_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 p_vLED_obuft_RNO_2_LC_11_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2833),
            .lcout(N_423_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ballX_RNICMG91_1_LC_11_7_0.C_ON=1'b0;
    defparam ballX_RNICMG91_1_LC_11_7_0.SEQ_MODE=4'b0000;
    defparam ballX_RNICMG91_1_LC_11_7_0.LUT_INIT=16'b1001000000001001;
    LogicCell40 ballX_RNICMG91_1_LC_11_7_0 (
            .in0(N__2812),
            .in1(N__3337),
            .in2(N__2791),
            .in3(N__3451),
            .lcout(p_hLED52_NE_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ballX_RNI38OK_0_LC_11_7_1.C_ON=1'b0;
    defparam ballX_RNI38OK_0_LC_11_7_1.SEQ_MODE=4'b0000;
    defparam ballX_RNI38OK_0_LC_11_7_1.LUT_INIT=16'b0011001111001100;
    LogicCell40 ballX_RNI38OK_0_LC_11_7_1 (
            .in0(_gnd_net_),
            .in1(N__2764),
            .in2(_gnd_net_),
            .in3(N__3230),
            .lcout(N_70_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ballX_RNIOC1J2_3_LC_11_8_4.C_ON=1'b0;
    defparam ballX_RNIOC1J2_3_LC_11_8_4.SEQ_MODE=4'b0000;
    defparam ballX_RNIOC1J2_3_LC_11_8_4.LUT_INIT=16'b0010000000000010;
    LogicCell40 ballX_RNIOC1J2_3_LC_11_8_4 (
            .in0(N__2746),
            .in1(N__2740),
            .in2(N__2734),
            .in3(N__3572),
            .lcout(p_hLED52),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam p_hLED_obuft_RNO_4_LC_11_8_5.C_ON=1'b0;
    defparam p_hLED_obuft_RNO_4_LC_11_8_5.SEQ_MODE=4'b0000;
    defparam p_hLED_obuft_RNO_4_LC_11_8_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 p_hLED_obuft_RNO_4_LC_11_8_5 (
            .in0(N__2914),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_410_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam p_hLED_cl_6_i_0_LC_11_9_0.C_ON=1'b0;
    defparam p_hLED_cl_6_i_0_LC_11_9_0.SEQ_MODE=4'b1000;
    defparam p_hLED_cl_6_i_0_LC_11_9_0.LUT_INIT=16'b1111111111111101;
    LogicCell40 p_hLED_cl_6_i_0_LC_11_9_0 (
            .in0(N__3486),
            .in1(N__3285),
            .in2(N__3409),
            .in3(N__3576),
            .lcout(p_hLED_cl_6_iZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3176),
            .ce(N__3136),
            .sr(_gnd_net_));
    defparam p_hLED_cl_4_i_0_LC_11_9_2.C_ON=1'b0;
    defparam p_hLED_cl_4_i_0_LC_11_9_2.SEQ_MODE=4'b1000;
    defparam p_hLED_cl_4_i_0_LC_11_9_2.LUT_INIT=16'b1111111111101111;
    LogicCell40 p_hLED_cl_4_i_0_LC_11_9_2 (
            .in0(N__3485),
            .in1(N__3284),
            .in2(N__3408),
            .in3(N__3575),
            .lcout(p_hLED_cl_4_iZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3176),
            .ce(N__3136),
            .sr(_gnd_net_));
    defparam p_hLED_cl_12_i_0_LC_11_9_6.C_ON=1'b0;
    defparam p_hLED_cl_12_i_0_LC_11_9_6.SEQ_MODE=4'b1000;
    defparam p_hLED_cl_12_i_0_LC_11_9_6.LUT_INIT=16'b1111101111111111;
    LogicCell40 p_hLED_cl_12_i_0_LC_11_9_6 (
            .in0(N__3484),
            .in1(N__3283),
            .in2(N__3407),
            .in3(N__3574),
            .lcout(p_hLED_cl_12_iZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3176),
            .ce(N__3136),
            .sr(_gnd_net_));
    defparam p_hLED_cl_8_i_0_LC_11_9_7.C_ON=1'b0;
    defparam p_hLED_cl_8_i_0_LC_11_9_7.SEQ_MODE=4'b1000;
    defparam p_hLED_cl_8_i_0_LC_11_9_7.LUT_INIT=16'b1110111111111111;
    LogicCell40 p_hLED_cl_8_i_0_LC_11_9_7 (
            .in0(N__3573),
            .in1(N__3380),
            .in2(N__3292),
            .in3(N__3487),
            .lcout(p_hLED_cl_8_iZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3176),
            .ce(N__3136),
            .sr(_gnd_net_));
    defparam p_vLED_obuft_RNO_6_LC_12_2_3.C_ON=1'b0;
    defparam p_vLED_obuft_RNO_6_LC_12_2_3.SEQ_MODE=4'b0000;
    defparam p_vLED_obuft_RNO_6_LC_12_2_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 p_vLED_obuft_RNO_6_LC_12_2_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2908),
            .lcout(N_427_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam p_vLED_obuft_RNO_5_LC_12_3_6.C_ON=1'b0;
    defparam p_vLED_obuft_RNO_5_LC_12_3_6.SEQ_MODE=4'b0000;
    defparam p_vLED_obuft_RNO_5_LC_12_3_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 p_vLED_obuft_RNO_5_LC_12_3_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2890),
            .lcout(N_426_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam p_hLED_obuft_RNO_8_LC_12_4_5.C_ON=1'b0;
    defparam p_hLED_obuft_RNO_8_LC_12_4_5.SEQ_MODE=4'b0000;
    defparam p_hLED_obuft_RNO_8_LC_12_4_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 p_hLED_obuft_RNO_8_LC_12_4_5 (
            .in0(N__2983),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_414_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam p_vLED_obuft_RNO_0_LC_12_5_3.C_ON=1'b0;
    defparam p_vLED_obuft_RNO_0_LC_12_5_3.SEQ_MODE=4'b0000;
    defparam p_vLED_obuft_RNO_0_LC_12_5_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 p_vLED_obuft_RNO_0_LC_12_5_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2860),
            .lcout(N_421_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_12_5_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_5_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_5_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam p_hLED_cl_7_i_0_LC_12_7_1.C_ON=1'b0;
    defparam p_hLED_cl_7_i_0_LC_12_7_1.SEQ_MODE=4'b1000;
    defparam p_hLED_cl_7_i_0_LC_12_7_1.LUT_INIT=16'b1111111111101110;
    LogicCell40 p_hLED_cl_7_i_0_LC_12_7_1 (
            .in0(N__3563),
            .in1(N__2974),
            .in2(_gnd_net_),
            .in3(N__3247),
            .lcout(p_hLED_cl_7_iZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3179),
            .ce(N__3131),
            .sr(_gnd_net_));
    defparam p_hLED_cl_i_0_LC_12_7_2.C_ON=1'b0;
    defparam p_hLED_cl_i_0_LC_12_7_2.SEQ_MODE=4'b1000;
    defparam p_hLED_cl_i_0_LC_12_7_2.LUT_INIT=16'b1111111011111111;
    LogicCell40 p_hLED_cl_i_0_LC_12_7_2 (
            .in0(N__3481),
            .in1(N__3242),
            .in2(N__3405),
            .in3(N__3567),
            .lcout(p_hLED_cl_iZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3179),
            .ce(N__3131),
            .sr(_gnd_net_));
    defparam p_hLED_cl_2_i_0_LC_12_7_3.C_ON=1'b0;
    defparam p_hLED_cl_2_i_0_LC_12_7_3.SEQ_MODE=4'b1000;
    defparam p_hLED_cl_2_i_0_LC_12_7_3.LUT_INIT=16'b1110111111111111;
    LogicCell40 p_hLED_cl_2_i_0_LC_12_7_3 (
            .in0(N__3564),
            .in1(N__3482),
            .in2(N__3406),
            .in3(N__3246),
            .lcout(p_hLED_cl_2_iZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3179),
            .ce(N__3131),
            .sr(_gnd_net_));
    defparam p_hLED_cl_1_i_0_LC_12_7_4.C_ON=1'b0;
    defparam p_hLED_cl_1_i_0_LC_12_7_4.SEQ_MODE=4'b1000;
    defparam p_hLED_cl_1_i_0_LC_12_7_4.LUT_INIT=16'b1111111110111011;
    LogicCell40 p_hLED_cl_1_i_0_LC_12_7_4 (
            .in0(N__2973),
            .in1(N__3243),
            .in2(_gnd_net_),
            .in3(N__3565),
            .lcout(p_hLED_cl_1_iZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3179),
            .ce(N__3131),
            .sr(_gnd_net_));
    defparam p_hLED_cl_14_i_0_LC_12_7_6.C_ON=1'b0;
    defparam p_hLED_cl_14_i_0_LC_12_7_6.SEQ_MODE=4'b1000;
    defparam p_hLED_cl_14_i_0_LC_12_7_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 p_hLED_cl_14_i_0_LC_12_7_6 (
            .in0(N__3480),
            .in1(N__3241),
            .in2(N__3404),
            .in3(N__3566),
            .lcout(p_hLED_cl_14_iZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3179),
            .ce(N__3131),
            .sr(_gnd_net_));
    defparam p_hLED_obuft_RNO_0_LC_12_8_0.C_ON=1'b0;
    defparam p_hLED_obuft_RNO_0_LC_12_8_0.SEQ_MODE=4'b0000;
    defparam p_hLED_obuft_RNO_0_LC_12_8_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 p_hLED_obuft_RNO_0_LC_12_8_0 (
            .in0(N__2959),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_406_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam p_hLED_obuft_RNO_2_LC_12_8_2.C_ON=1'b0;
    defparam p_hLED_obuft_RNO_2_LC_12_8_2.SEQ_MODE=4'b0000;
    defparam p_hLED_obuft_RNO_2_LC_12_8_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 p_hLED_obuft_RNO_2_LC_12_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2947),
            .lcout(N_408_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam p_hLED_obuft_RNO_1_LC_12_8_4.C_ON=1'b0;
    defparam p_hLED_obuft_RNO_1_LC_12_8_4.SEQ_MODE=4'b0000;
    defparam p_hLED_obuft_RNO_1_LC_12_8_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 p_hLED_obuft_RNO_1_LC_12_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3592),
            .lcout(N_407_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam p_hLED_obuft_RNO_3_LC_12_8_7.C_ON=1'b0;
    defparam p_hLED_obuft_RNO_3_LC_12_8_7.SEQ_MODE=4'b0000;
    defparam p_hLED_obuft_RNO_3_LC_12_8_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 p_hLED_obuft_RNO_3_LC_12_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3604),
            .lcout(N_409_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam p_hLED_cl_10_i_0_LC_12_9_0.C_ON=1'b0;
    defparam p_hLED_cl_10_i_0_LC_12_9_0.SEQ_MODE=4'b1000;
    defparam p_hLED_cl_10_i_0_LC_12_9_0.LUT_INIT=16'b1011111111111111;
    LogicCell40 p_hLED_cl_10_i_0_LC_12_9_0 (
            .in0(N__3488),
            .in1(N__3584),
            .in2(N__3289),
            .in3(N__3399),
            .lcout(p_hLED_cl_10_iZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3180),
            .ce(N__3135),
            .sr(_gnd_net_));
    defparam p_hLED_cl_9_i_0_LC_12_9_1.C_ON=1'b0;
    defparam p_hLED_cl_9_i_0_LC_12_9_1.SEQ_MODE=4'b1000;
    defparam p_hLED_cl_9_i_0_LC_12_9_1.LUT_INIT=16'b1111111111110111;
    LogicCell40 p_hLED_cl_9_i_0_LC_12_9_1 (
            .in0(N__3582),
            .in1(N__3493),
            .in2(N__3412),
            .in3(N__3282),
            .lcout(p_hLED_cl_9_iZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3180),
            .ce(N__3135),
            .sr(_gnd_net_));
    defparam p_hLED_cl_3_i_0_LC_12_9_3.C_ON=1'b0;
    defparam p_hLED_cl_3_i_0_LC_12_9_3.SEQ_MODE=4'b1000;
    defparam p_hLED_cl_3_i_0_LC_12_9_3.LUT_INIT=16'b1111111011111111;
    LogicCell40 p_hLED_cl_3_i_0_LC_12_9_3 (
            .in0(N__3581),
            .in1(N__3492),
            .in2(N__3411),
            .in3(N__3281),
            .lcout(p_hLED_cl_3_iZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3180),
            .ce(N__3135),
            .sr(_gnd_net_));
    defparam p_hLED_cl_11_i_0_LC_12_9_4.C_ON=1'b0;
    defparam p_hLED_cl_11_i_0_LC_12_9_4.SEQ_MODE=4'b1000;
    defparam p_hLED_cl_11_i_0_LC_12_9_4.LUT_INIT=16'b1111011111111111;
    LogicCell40 p_hLED_cl_11_i_0_LC_12_9_4 (
            .in0(N__3489),
            .in1(N__3583),
            .in2(N__3291),
            .in3(N__3401),
            .lcout(p_hLED_cl_11_iZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3180),
            .ce(N__3135),
            .sr(_gnd_net_));
    defparam p_hLED_cl_5_i_0_LC_12_9_6.C_ON=1'b0;
    defparam p_hLED_cl_5_i_0_LC_12_9_6.SEQ_MODE=4'b1000;
    defparam p_hLED_cl_5_i_0_LC_12_9_6.LUT_INIT=16'b1111111101111111;
    LogicCell40 p_hLED_cl_5_i_0_LC_12_9_6 (
            .in0(N__3490),
            .in1(N__3585),
            .in2(N__3290),
            .in3(N__3400),
            .lcout(p_hLED_cl_5_iZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3180),
            .ce(N__3135),
            .sr(_gnd_net_));
    defparam p_hLED_cl_13_i_0_LC_12_9_7.C_ON=1'b0;
    defparam p_hLED_cl_13_i_0_LC_12_9_7.SEQ_MODE=4'b1000;
    defparam p_hLED_cl_13_i_0_LC_12_9_7.LUT_INIT=16'b1111111111011111;
    LogicCell40 p_hLED_cl_13_i_0_LC_12_9_7 (
            .in0(N__3580),
            .in1(N__3491),
            .in2(N__3410),
            .in3(N__3280),
            .lcout(p_hLED_cl_13_iZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3180),
            .ce(N__3135),
            .sr(_gnd_net_));
    defparam p_hLED_obuft_RNO_10_LC_12_10_4.C_ON=1'b0;
    defparam p_hLED_obuft_RNO_10_LC_12_10_4.SEQ_MODE=4'b0000;
    defparam p_hLED_obuft_RNO_10_LC_12_10_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 p_hLED_obuft_RNO_10_LC_12_10_4 (
            .in0(N__3103),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_416_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam p_hLED_obuft_RNO_5_LC_12_10_5.C_ON=1'b0;
    defparam p_hLED_obuft_RNO_5_LC_12_10_5.SEQ_MODE=4'b0000;
    defparam p_hLED_obuft_RNO_5_LC_12_10_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 p_hLED_obuft_RNO_5_LC_12_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3085),
            .lcout(N_411_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam p_hLED_obuft_RNO_11_LC_12_10_7.C_ON=1'b0;
    defparam p_hLED_obuft_RNO_11_LC_12_10_7.SEQ_MODE=4'b0000;
    defparam p_hLED_obuft_RNO_11_LC_12_10_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 p_hLED_obuft_RNO_11_LC_12_10_7 (
            .in0(N__3721),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_417_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam p_hLED_obuft_RNO_12_LC_12_11_1.C_ON=1'b0;
    defparam p_hLED_obuft_RNO_12_LC_12_11_1.SEQ_MODE=4'b0000;
    defparam p_hLED_obuft_RNO_12_LC_12_11_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 p_hLED_obuft_RNO_12_LC_12_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3700),
            .lcout(N_418_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam p_hLED_obuft_RNO_7_LC_12_12_4.C_ON=1'b0;
    defparam p_hLED_obuft_RNO_7_LC_12_12_4.SEQ_MODE=4'b0000;
    defparam p_hLED_obuft_RNO_7_LC_12_12_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 p_hLED_obuft_RNO_7_LC_12_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3676),
            .lcout(N_413_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam p_hLED_obuft_RNO_14_LC_12_13_0.C_ON=1'b0;
    defparam p_hLED_obuft_RNO_14_LC_12_13_0.SEQ_MODE=4'b0000;
    defparam p_hLED_obuft_RNO_14_LC_12_13_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 p_hLED_obuft_RNO_14_LC_12_13_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3658),
            .lcout(N_420_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam p_hLED_obuft_RNO_9_LC_12_13_5.C_ON=1'b0;
    defparam p_hLED_obuft_RNO_9_LC_12_13_5.SEQ_MODE=4'b0000;
    defparam p_hLED_obuft_RNO_9_LC_12_13_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 p_hLED_obuft_RNO_9_LC_12_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3637),
            .lcout(N_415_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam p_hLED_obuft_RNO_13_LC_12_15_0.C_ON=1'b0;
    defparam p_hLED_obuft_RNO_13_LC_12_15_0.SEQ_MODE=4'b0000;
    defparam p_hLED_obuft_RNO_13_LC_12_15_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 p_hLED_obuft_RNO_13_LC_12_15_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3619),
            .lcout(N_419_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // top
