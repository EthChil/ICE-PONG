-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Dec 13 2020 21:22:15

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    p_hLED : out std_logic_vector(14 downto 0);
    p_vLED : out std_logic_vector(9 downto 0);
    p_dwnBtn : in std_logic;
    p_upBtn : in std_logic;
    p_clk12 : in std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__3967\ : std_logic;
signal \N__3966\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3956\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3946\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3938\ : std_logic;
signal \N__3937\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3929\ : std_logic;
signal \N__3928\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3919\ : std_logic;
signal \N__3918\ : std_logic;
signal \N__3911\ : std_logic;
signal \N__3910\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3901\ : std_logic;
signal \N__3900\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3892\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3874\ : std_logic;
signal \N__3873\ : std_logic;
signal \N__3866\ : std_logic;
signal \N__3865\ : std_logic;
signal \N__3864\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3856\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3847\ : std_logic;
signal \N__3846\ : std_logic;
signal \N__3839\ : std_logic;
signal \N__3838\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3829\ : std_logic;
signal \N__3828\ : std_logic;
signal \N__3821\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3811\ : std_logic;
signal \N__3810\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3802\ : std_logic;
signal \N__3801\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3793\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3785\ : std_logic;
signal \N__3784\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3776\ : std_logic;
signal \N__3775\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3767\ : std_logic;
signal \N__3766\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3758\ : std_logic;
signal \N__3757\ : std_logic;
signal \N__3756\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3748\ : std_logic;
signal \N__3747\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3738\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3718\ : std_logic;
signal \N__3715\ : std_logic;
signal \N__3712\ : std_logic;
signal \N__3709\ : std_logic;
signal \N__3706\ : std_logic;
signal \N__3703\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3694\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3688\ : std_logic;
signal \N__3685\ : std_logic;
signal \N__3682\ : std_logic;
signal \N__3679\ : std_logic;
signal \N__3676\ : std_logic;
signal \N__3673\ : std_logic;
signal \N__3670\ : std_logic;
signal \N__3667\ : std_logic;
signal \N__3664\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3655\ : std_logic;
signal \N__3652\ : std_logic;
signal \N__3649\ : std_logic;
signal \N__3646\ : std_logic;
signal \N__3643\ : std_logic;
signal \N__3640\ : std_logic;
signal \N__3637\ : std_logic;
signal \N__3634\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3625\ : std_logic;
signal \N__3622\ : std_logic;
signal \N__3619\ : std_logic;
signal \N__3616\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3607\ : std_logic;
signal \N__3604\ : std_logic;
signal \N__3601\ : std_logic;
signal \N__3598\ : std_logic;
signal \N__3595\ : std_logic;
signal \N__3592\ : std_logic;
signal \N__3589\ : std_logic;
signal \N__3586\ : std_logic;
signal \N__3585\ : std_logic;
signal \N__3584\ : std_logic;
signal \N__3583\ : std_logic;
signal \N__3582\ : std_logic;
signal \N__3581\ : std_logic;
signal \N__3580\ : std_logic;
signal \N__3577\ : std_logic;
signal \N__3576\ : std_logic;
signal \N__3575\ : std_logic;
signal \N__3574\ : std_logic;
signal \N__3573\ : std_logic;
signal \N__3572\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3570\ : std_logic;
signal \N__3569\ : std_logic;
signal \N__3568\ : std_logic;
signal \N__3567\ : std_logic;
signal \N__3566\ : std_logic;
signal \N__3565\ : std_logic;
signal \N__3564\ : std_logic;
signal \N__3563\ : std_logic;
signal \N__3550\ : std_logic;
signal \N__3547\ : std_logic;
signal \N__3538\ : std_logic;
signal \N__3535\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3515\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3509\ : std_logic;
signal \N__3504\ : std_logic;
signal \N__3493\ : std_logic;
signal \N__3492\ : std_logic;
signal \N__3491\ : std_logic;
signal \N__3490\ : std_logic;
signal \N__3489\ : std_logic;
signal \N__3488\ : std_logic;
signal \N__3487\ : std_logic;
signal \N__3486\ : std_logic;
signal \N__3485\ : std_logic;
signal \N__3484\ : std_logic;
signal \N__3483\ : std_logic;
signal \N__3482\ : std_logic;
signal \N__3481\ : std_logic;
signal \N__3480\ : std_logic;
signal \N__3467\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3457\ : std_logic;
signal \N__3456\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3452\ : std_logic;
signal \N__3451\ : std_logic;
signal \N__3444\ : std_logic;
signal \N__3441\ : std_logic;
signal \N__3438\ : std_logic;
signal \N__3431\ : std_logic;
signal \N__3428\ : std_logic;
signal \N__3425\ : std_logic;
signal \N__3412\ : std_logic;
signal \N__3411\ : std_logic;
signal \N__3410\ : std_logic;
signal \N__3409\ : std_logic;
signal \N__3408\ : std_logic;
signal \N__3407\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3404\ : std_logic;
signal \N__3403\ : std_logic;
signal \N__3402\ : std_logic;
signal \N__3401\ : std_logic;
signal \N__3400\ : std_logic;
signal \N__3399\ : std_logic;
signal \N__3396\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3390\ : std_logic;
signal \N__3387\ : std_logic;
signal \N__3384\ : std_logic;
signal \N__3381\ : std_logic;
signal \N__3380\ : std_logic;
signal \N__3379\ : std_logic;
signal \N__3376\ : std_logic;
signal \N__3373\ : std_logic;
signal \N__3370\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3342\ : std_logic;
signal \N__3341\ : std_logic;
signal \N__3338\ : std_logic;
signal \N__3337\ : std_logic;
signal \N__3334\ : std_logic;
signal \N__3329\ : std_logic;
signal \N__3324\ : std_logic;
signal \N__3321\ : std_logic;
signal \N__3318\ : std_logic;
signal \N__3315\ : std_logic;
signal \N__3312\ : std_logic;
signal \N__3309\ : std_logic;
signal \N__3292\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3290\ : std_logic;
signal \N__3289\ : std_logic;
signal \N__3286\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3284\ : std_logic;
signal \N__3283\ : std_logic;
signal \N__3282\ : std_logic;
signal \N__3281\ : std_logic;
signal \N__3280\ : std_logic;
signal \N__3277\ : std_logic;
signal \N__3274\ : std_logic;
signal \N__3271\ : std_logic;
signal \N__3262\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3248\ : std_logic;
signal \N__3247\ : std_logic;
signal \N__3246\ : std_logic;
signal \N__3245\ : std_logic;
signal \N__3244\ : std_logic;
signal \N__3243\ : std_logic;
signal \N__3242\ : std_logic;
signal \N__3241\ : std_logic;
signal \N__3240\ : std_logic;
signal \N__3239\ : std_logic;
signal \N__3234\ : std_logic;
signal \N__3231\ : std_logic;
signal \N__3230\ : std_logic;
signal \N__3225\ : std_logic;
signal \N__3220\ : std_logic;
signal \N__3213\ : std_logic;
signal \N__3210\ : std_logic;
signal \N__3207\ : std_logic;
signal \N__3204\ : std_logic;
signal \N__3201\ : std_logic;
signal \N__3198\ : std_logic;
signal \N__3181\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3179\ : std_logic;
signal \N__3178\ : std_logic;
signal \N__3177\ : std_logic;
signal \N__3176\ : std_logic;
signal \N__3175\ : std_logic;
signal \N__3174\ : std_logic;
signal \N__3173\ : std_logic;
signal \N__3172\ : std_logic;
signal \N__3171\ : std_logic;
signal \N__3170\ : std_logic;
signal \N__3169\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3135\ : std_logic;
signal \N__3132\ : std_logic;
signal \N__3131\ : std_logic;
signal \N__3128\ : std_logic;
signal \N__3125\ : std_logic;
signal \N__3122\ : std_logic;
signal \N__3119\ : std_logic;
signal \N__3114\ : std_logic;
signal \N__3109\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3103\ : std_logic;
signal \N__3100\ : std_logic;
signal \N__3097\ : std_logic;
signal \N__3094\ : std_logic;
signal \N__3091\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3085\ : std_logic;
signal \N__3082\ : std_logic;
signal \N__3079\ : std_logic;
signal \N__3076\ : std_logic;
signal \N__3073\ : std_logic;
signal \N__3072\ : std_logic;
signal \N__3071\ : std_logic;
signal \N__3070\ : std_logic;
signal \N__3067\ : std_logic;
signal \N__3064\ : std_logic;
signal \N__3063\ : std_logic;
signal \N__3062\ : std_logic;
signal \N__3059\ : std_logic;
signal \N__3056\ : std_logic;
signal \N__3051\ : std_logic;
signal \N__3048\ : std_logic;
signal \N__3045\ : std_logic;
signal \N__3038\ : std_logic;
signal \N__3035\ : std_logic;
signal \N__3032\ : std_logic;
signal \N__3031\ : std_logic;
signal \N__3030\ : std_logic;
signal \N__3029\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3020\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3014\ : std_logic;
signal \N__3011\ : std_logic;
signal \N__3008\ : std_logic;
signal \N__2995\ : std_logic;
signal \N__2992\ : std_logic;
signal \N__2989\ : std_logic;
signal \N__2986\ : std_logic;
signal \N__2983\ : std_logic;
signal \N__2980\ : std_logic;
signal \N__2977\ : std_logic;
signal \N__2974\ : std_logic;
signal \N__2973\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2967\ : std_logic;
signal \N__2964\ : std_logic;
signal \N__2959\ : std_logic;
signal \N__2956\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2950\ : std_logic;
signal \N__2947\ : std_logic;
signal \N__2944\ : std_logic;
signal \N__2941\ : std_logic;
signal \N__2938\ : std_logic;
signal \N__2935\ : std_logic;
signal \N__2932\ : std_logic;
signal \N__2929\ : std_logic;
signal \N__2926\ : std_logic;
signal \N__2923\ : std_logic;
signal \N__2920\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2914\ : std_logic;
signal \N__2911\ : std_logic;
signal \N__2908\ : std_logic;
signal \N__2905\ : std_logic;
signal \N__2902\ : std_logic;
signal \N__2899\ : std_logic;
signal \N__2896\ : std_logic;
signal \N__2893\ : std_logic;
signal \N__2890\ : std_logic;
signal \N__2887\ : std_logic;
signal \N__2884\ : std_logic;
signal \N__2881\ : std_logic;
signal \N__2878\ : std_logic;
signal \N__2875\ : std_logic;
signal \N__2872\ : std_logic;
signal \N__2869\ : std_logic;
signal \N__2866\ : std_logic;
signal \N__2863\ : std_logic;
signal \N__2860\ : std_logic;
signal \N__2857\ : std_logic;
signal \N__2854\ : std_logic;
signal \N__2851\ : std_logic;
signal \N__2848\ : std_logic;
signal \N__2845\ : std_logic;
signal \N__2842\ : std_logic;
signal \N__2839\ : std_logic;
signal \N__2836\ : std_logic;
signal \N__2833\ : std_logic;
signal \N__2830\ : std_logic;
signal \N__2827\ : std_logic;
signal \N__2824\ : std_logic;
signal \N__2821\ : std_logic;
signal \N__2818\ : std_logic;
signal \N__2815\ : std_logic;
signal \N__2812\ : std_logic;
signal \N__2811\ : std_logic;
signal \N__2810\ : std_logic;
signal \N__2807\ : std_logic;
signal \N__2804\ : std_logic;
signal \N__2801\ : std_logic;
signal \N__2798\ : std_logic;
signal \N__2791\ : std_logic;
signal \N__2790\ : std_logic;
signal \N__2787\ : std_logic;
signal \N__2786\ : std_logic;
signal \N__2783\ : std_logic;
signal \N__2780\ : std_logic;
signal \N__2777\ : std_logic;
signal \N__2774\ : std_logic;
signal \N__2771\ : std_logic;
signal \N__2764\ : std_logic;
signal \N__2763\ : std_logic;
signal \N__2762\ : std_logic;
signal \N__2759\ : std_logic;
signal \N__2754\ : std_logic;
signal \N__2751\ : std_logic;
signal \N__2746\ : std_logic;
signal \N__2743\ : std_logic;
signal \N__2740\ : std_logic;
signal \N__2737\ : std_logic;
signal \N__2734\ : std_logic;
signal \N__2731\ : std_logic;
signal \N__2728\ : std_logic;
signal \N__2727\ : std_logic;
signal \N__2726\ : std_logic;
signal \N__2723\ : std_logic;
signal \N__2718\ : std_logic;
signal \N__2715\ : std_logic;
signal \N__2710\ : std_logic;
signal \N__2709\ : std_logic;
signal \N__2706\ : std_logic;
signal \N__2703\ : std_logic;
signal \N__2700\ : std_logic;
signal \N__2695\ : std_logic;
signal \N__2692\ : std_logic;
signal \N__2689\ : std_logic;
signal \N__2688\ : std_logic;
signal \N__2685\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2679\ : std_logic;
signal \N__2674\ : std_logic;
signal \N__2671\ : std_logic;
signal \N__2668\ : std_logic;
signal \N__2667\ : std_logic;
signal \N__2664\ : std_logic;
signal \N__2661\ : std_logic;
signal \N__2658\ : std_logic;
signal \N__2653\ : std_logic;
signal \N__2650\ : std_logic;
signal \N__2647\ : std_logic;
signal \N__2646\ : std_logic;
signal \N__2643\ : std_logic;
signal \N__2640\ : std_logic;
signal \N__2637\ : std_logic;
signal \N__2632\ : std_logic;
signal \N__2629\ : std_logic;
signal \N__2626\ : std_logic;
signal \N__2623\ : std_logic;
signal \N__2620\ : std_logic;
signal \N__2617\ : std_logic;
signal \N__2614\ : std_logic;
signal \N__2611\ : std_logic;
signal \N__2608\ : std_logic;
signal \N__2605\ : std_logic;
signal \N__2602\ : std_logic;
signal \N__2599\ : std_logic;
signal \N__2596\ : std_logic;
signal \N__2593\ : std_logic;
signal \N__2590\ : std_logic;
signal \N__2587\ : std_logic;
signal \N__2584\ : std_logic;
signal \N__2581\ : std_logic;
signal \N__2578\ : std_logic;
signal \N__2575\ : std_logic;
signal \N__2572\ : std_logic;
signal \N__2569\ : std_logic;
signal \N__2566\ : std_logic;
signal \N__2563\ : std_logic;
signal \N__2560\ : std_logic;
signal \N__2557\ : std_logic;
signal \N__2554\ : std_logic;
signal \N__2551\ : std_logic;
signal \N__2548\ : std_logic;
signal \N__2545\ : std_logic;
signal \N__2542\ : std_logic;
signal \N__2539\ : std_logic;
signal \N__2538\ : std_logic;
signal \N__2535\ : std_logic;
signal \N__2532\ : std_logic;
signal \N__2529\ : std_logic;
signal \N__2524\ : std_logic;
signal \N__2521\ : std_logic;
signal \N__2518\ : std_logic;
signal \N__2517\ : std_logic;
signal \N__2514\ : std_logic;
signal \N__2511\ : std_logic;
signal \N__2506\ : std_logic;
signal \N__2503\ : std_logic;
signal \N__2502\ : std_logic;
signal \N__2499\ : std_logic;
signal \N__2496\ : std_logic;
signal \N__2493\ : std_logic;
signal \N__2488\ : std_logic;
signal \N__2485\ : std_logic;
signal \N__2484\ : std_logic;
signal \N__2481\ : std_logic;
signal \N__2478\ : std_logic;
signal \N__2473\ : std_logic;
signal \N__2470\ : std_logic;
signal \N__2469\ : std_logic;
signal \N__2466\ : std_logic;
signal \N__2463\ : std_logic;
signal \N__2458\ : std_logic;
signal \N__2455\ : std_logic;
signal \N__2454\ : std_logic;
signal \N__2451\ : std_logic;
signal \N__2448\ : std_logic;
signal \N__2443\ : std_logic;
signal \N__2440\ : std_logic;
signal \N__2439\ : std_logic;
signal \N__2436\ : std_logic;
signal \N__2433\ : std_logic;
signal \N__2428\ : std_logic;
signal \N__2425\ : std_logic;
signal \N__2424\ : std_logic;
signal \N__2421\ : std_logic;
signal \N__2418\ : std_logic;
signal \N__2415\ : std_logic;
signal \N__2410\ : std_logic;
signal \N__2407\ : std_logic;
signal \N__2406\ : std_logic;
signal \N__2405\ : std_logic;
signal \N__2404\ : std_logic;
signal \N__2401\ : std_logic;
signal \N__2398\ : std_logic;
signal \N__2395\ : std_logic;
signal \N__2392\ : std_logic;
signal \N__2383\ : std_logic;
signal \N__2380\ : std_logic;
signal \N__2377\ : std_logic;
signal \N__2376\ : std_logic;
signal \N__2373\ : std_logic;
signal \N__2370\ : std_logic;
signal \N__2365\ : std_logic;
signal \N__2364\ : std_logic;
signal \N__2363\ : std_logic;
signal \N__2362\ : std_logic;
signal \N__2361\ : std_logic;
signal \N__2360\ : std_logic;
signal \N__2359\ : std_logic;
signal \N__2346\ : std_logic;
signal \N__2345\ : std_logic;
signal \N__2344\ : std_logic;
signal \N__2343\ : std_logic;
signal \N__2340\ : std_logic;
signal \N__2339\ : std_logic;
signal \N__2338\ : std_logic;
signal \N__2335\ : std_logic;
signal \N__2328\ : std_logic;
signal \N__2325\ : std_logic;
signal \N__2320\ : std_logic;
signal \N__2311\ : std_logic;
signal \N__2310\ : std_logic;
signal \N__2307\ : std_logic;
signal \N__2304\ : std_logic;
signal \N__2299\ : std_logic;
signal \N__2296\ : std_logic;
signal \N__2293\ : std_logic;
signal \N__2292\ : std_logic;
signal \N__2289\ : std_logic;
signal \N__2286\ : std_logic;
signal \N__2283\ : std_logic;
signal \N__2278\ : std_logic;
signal \N__2275\ : std_logic;
signal \N__2274\ : std_logic;
signal \N__2271\ : std_logic;
signal \N__2268\ : std_logic;
signal \N__2263\ : std_logic;
signal \N__2260\ : std_logic;
signal \N__2259\ : std_logic;
signal \N__2256\ : std_logic;
signal \N__2253\ : std_logic;
signal \N__2248\ : std_logic;
signal \N__2245\ : std_logic;
signal \N__2244\ : std_logic;
signal \N__2241\ : std_logic;
signal \N__2238\ : std_logic;
signal \N__2233\ : std_logic;
signal \N__2230\ : std_logic;
signal \N__2229\ : std_logic;
signal \N__2226\ : std_logic;
signal \N__2223\ : std_logic;
signal \N__2218\ : std_logic;
signal \N__2215\ : std_logic;
signal \N__2214\ : std_logic;
signal \N__2211\ : std_logic;
signal \N__2208\ : std_logic;
signal \N__2205\ : std_logic;
signal \N__2200\ : std_logic;
signal \N__2197\ : std_logic;
signal \N__2194\ : std_logic;
signal \N__2191\ : std_logic;
signal \N__2188\ : std_logic;
signal \N__2185\ : std_logic;
signal \N__2182\ : std_logic;
signal \N__2179\ : std_logic;
signal \N__2178\ : std_logic;
signal \N__2175\ : std_logic;
signal \N__2172\ : std_logic;
signal \N__2169\ : std_logic;
signal \N__2166\ : std_logic;
signal \N__2161\ : std_logic;
signal \N__2160\ : std_logic;
signal \N__2159\ : std_logic;
signal \N__2158\ : std_logic;
signal \N__2157\ : std_logic;
signal \N__2156\ : std_logic;
signal \N__2155\ : std_logic;
signal \N__2154\ : std_logic;
signal \N__2141\ : std_logic;
signal \N__2140\ : std_logic;
signal \N__2139\ : std_logic;
signal \N__2138\ : std_logic;
signal \N__2135\ : std_logic;
signal \N__2134\ : std_logic;
signal \N__2131\ : std_logic;
signal \N__2128\ : std_logic;
signal \N__2121\ : std_logic;
signal \N__2116\ : std_logic;
signal \N__2113\ : std_logic;
signal \N__2104\ : std_logic;
signal \N__2103\ : std_logic;
signal \N__2102\ : std_logic;
signal \N__2101\ : std_logic;
signal \N__2100\ : std_logic;
signal \N__2097\ : std_logic;
signal \N__2094\ : std_logic;
signal \N__2091\ : std_logic;
signal \N__2090\ : std_logic;
signal \N__2089\ : std_logic;
signal \N__2088\ : std_logic;
signal \N__2085\ : std_logic;
signal \N__2082\ : std_logic;
signal \N__2081\ : std_logic;
signal \N__2068\ : std_logic;
signal \N__2067\ : std_logic;
signal \N__2066\ : std_logic;
signal \N__2065\ : std_logic;
signal \N__2058\ : std_logic;
signal \N__2055\ : std_logic;
signal \N__2052\ : std_logic;
signal \N__2049\ : std_logic;
signal \N__2046\ : std_logic;
signal \N__2035\ : std_logic;
signal \N__2034\ : std_logic;
signal \N__2033\ : std_logic;
signal \N__2032\ : std_logic;
signal \N__2031\ : std_logic;
signal \N__2030\ : std_logic;
signal \N__2027\ : std_logic;
signal \N__2024\ : std_logic;
signal \N__2021\ : std_logic;
signal \N__2020\ : std_logic;
signal \N__2019\ : std_logic;
signal \N__2006\ : std_logic;
signal \N__2005\ : std_logic;
signal \N__2004\ : std_logic;
signal \N__2001\ : std_logic;
signal \N__2000\ : std_logic;
signal \N__1999\ : std_logic;
signal \N__1996\ : std_logic;
signal \N__1993\ : std_logic;
signal \N__1986\ : std_logic;
signal \N__1983\ : std_logic;
signal \N__1980\ : std_logic;
signal \N__1977\ : std_logic;
signal \N__1966\ : std_logic;
signal \N__1963\ : std_logic;
signal \N__1960\ : std_logic;
signal \N__1957\ : std_logic;
signal \N__1954\ : std_logic;
signal \N__1951\ : std_logic;
signal \N__1948\ : std_logic;
signal \N__1945\ : std_logic;
signal \N__1942\ : std_logic;
signal \N__1939\ : std_logic;
signal \N__1938\ : std_logic;
signal \N__1937\ : std_logic;
signal \N__1936\ : std_logic;
signal \N__1933\ : std_logic;
signal \N__1932\ : std_logic;
signal \N__1931\ : std_logic;
signal \N__1928\ : std_logic;
signal \N__1927\ : std_logic;
signal \N__1926\ : std_logic;
signal \N__1925\ : std_logic;
signal \N__1922\ : std_logic;
signal \N__1921\ : std_logic;
signal \N__1918\ : std_logic;
signal \N__1913\ : std_logic;
signal \N__1904\ : std_logic;
signal \N__1897\ : std_logic;
signal \N__1888\ : std_logic;
signal \N__1885\ : std_logic;
signal \N__1882\ : std_logic;
signal \N__1879\ : std_logic;
signal \N__1876\ : std_logic;
signal \N__1873\ : std_logic;
signal \N__1870\ : std_logic;
signal \N__1867\ : std_logic;
signal \N__1864\ : std_logic;
signal \N__1861\ : std_logic;
signal \N__1858\ : std_logic;
signal \N__1855\ : std_logic;
signal \N__1852\ : std_logic;
signal \N__1849\ : std_logic;
signal \N__1848\ : std_logic;
signal \N__1847\ : std_logic;
signal \N__1844\ : std_logic;
signal \N__1839\ : std_logic;
signal \N__1834\ : std_logic;
signal \N__1831\ : std_logic;
signal \N__1830\ : std_logic;
signal \N__1829\ : std_logic;
signal \N__1826\ : std_logic;
signal \N__1823\ : std_logic;
signal \N__1820\ : std_logic;
signal \N__1813\ : std_logic;
signal \N__1810\ : std_logic;
signal \N__1809\ : std_logic;
signal \N__1808\ : std_logic;
signal \N__1807\ : std_logic;
signal \N__1806\ : std_logic;
signal \N__1803\ : std_logic;
signal \N__1798\ : std_logic;
signal \N__1793\ : std_logic;
signal \N__1786\ : std_logic;
signal \N__1785\ : std_logic;
signal \N__1782\ : std_logic;
signal \N__1781\ : std_logic;
signal \N__1778\ : std_logic;
signal \N__1773\ : std_logic;
signal \N__1768\ : std_logic;
signal \N__1767\ : std_logic;
signal \N__1764\ : std_logic;
signal \N__1763\ : std_logic;
signal \N__1760\ : std_logic;
signal \N__1757\ : std_logic;
signal \N__1752\ : std_logic;
signal \N__1747\ : std_logic;
signal \N__1744\ : std_logic;
signal \N__1741\ : std_logic;
signal \N__1738\ : std_logic;
signal \N__1735\ : std_logic;
signal \N__1732\ : std_logic;
signal \N__1729\ : std_logic;
signal \N__1726\ : std_logic;
signal \N__1723\ : std_logic;
signal \N__1720\ : std_logic;
signal \N__1717\ : std_logic;
signal \N__1716\ : std_logic;
signal \N__1715\ : std_logic;
signal \N__1714\ : std_logic;
signal \N__1713\ : std_logic;
signal \N__1702\ : std_logic;
signal \N__1699\ : std_logic;
signal \N__1696\ : std_logic;
signal \N__1693\ : std_logic;
signal \N__1690\ : std_logic;
signal \N__1687\ : std_logic;
signal \N__1684\ : std_logic;
signal \N__1681\ : std_logic;
signal \N__1678\ : std_logic;
signal \N__1675\ : std_logic;
signal \N__1672\ : std_logic;
signal \N__1669\ : std_logic;
signal \N__1666\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \bfn_7_6_0_\ : std_logic;
signal \un1_ballY_4_cry_0\ : std_logic;
signal \un1_ballY_4_cry_1\ : std_logic;
signal \un1_ballY_4_cry_2\ : std_logic;
signal \ballYVel_RNIGOGN4_0Z0Z_0\ : std_logic;
signal \ballYVel_RNIGOGN4Z0Z_0\ : std_logic;
signal \bfn_7_7_0_\ : std_logic;
signal \un1_ballX_3_cry_0\ : std_logic;
signal \un1_ballX_3_cry_1\ : std_logic;
signal \un1_ballX_3_cry_2\ : std_logic;
signal \ballXVel_s_1_0_0_cascade_\ : std_logic;
signal \ballXVel_RNIFI1J4_0Z0Z_0\ : std_logic;
signal \ballXVelZ0Z_0\ : std_logic;
signal \ballXVel_RNIFI1J4Z0Z_0\ : std_logic;
signal \N_67_i\ : std_logic;
signal \bfn_8_6_0_\ : std_logic;
signal \un1_vIndex_2_cry_0\ : std_logic;
signal \un1_vIndex_2_cry_1\ : std_logic;
signal \un1_vIndex_2_cry_2\ : std_logic;
signal \ballYZ0Z_0\ : std_logic;
signal \ballYZ0Z_1\ : std_logic;
signal \ballYVel_s_1_0_0_cascade_\ : std_logic;
signal \ballYVelZ0Z_0\ : std_logic;
signal \ballYZ0Z_2\ : std_logic;
signal \ballYZ0Z_3\ : std_logic;
signal \p_vLED37_NE_0\ : std_logic;
signal \ballXVel12_10_cascade_\ : std_logic;
signal \ballXVel12_12\ : std_logic;
signal \ballXVel12_14_cascade_\ : std_logic;
signal \ballXVel12_11\ : std_logic;
signal \ballXVel12\ : std_logic;
signal \ballXVel12_13\ : std_logic;
signal \N_430_i\ : std_logic;
signal \N_428_i\ : std_logic;
signal \p_vLED_cl_2_iZ0Z_0\ : std_logic;
signal \p_vLED_cl_9_iZ0Z_0\ : std_logic;
signal \p_vLED37\ : std_logic;
signal \vIndexZ0Z_2\ : std_logic;
signal \vIndexZ0Z_1\ : std_logic;
signal \vIndexZ0Z_3\ : std_logic;
signal \N_76_cascade_\ : std_logic;
signal \N_57_i\ : std_logic;
signal \p_vLED33\ : std_logic;
signal \N_57_i_cascade_\ : std_logic;
signal \N_76\ : std_logic;
signal \vIndexZ0Z_0\ : std_logic;
signal \ctrZ0Z_0\ : std_logic;
signal \bfn_9_7_0_\ : std_logic;
signal \ctrZ0Z_1\ : std_logic;
signal ctr_cry_0 : std_logic;
signal \ctrZ0Z_2\ : std_logic;
signal ctr_cry_1 : std_logic;
signal \ctrZ0Z_3\ : std_logic;
signal ctr_cry_2 : std_logic;
signal \ctrZ0Z_4\ : std_logic;
signal ctr_cry_3 : std_logic;
signal \ctrZ0Z_5\ : std_logic;
signal ctr_cry_4 : std_logic;
signal \ctrZ0Z_6\ : std_logic;
signal ctr_cry_5 : std_logic;
signal \ctrZ0Z_7\ : std_logic;
signal ctr_cry_6 : std_logic;
signal ctr_cry_7 : std_logic;
signal \ctrZ0Z_8\ : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \ctrZ0Z_9\ : std_logic;
signal ctr_cry_8 : std_logic;
signal \ctrZ0Z_10\ : std_logic;
signal ctr_cry_9 : std_logic;
signal \ctrZ0Z_11\ : std_logic;
signal ctr_cry_10 : std_logic;
signal \ctrZ0Z_12\ : std_logic;
signal ctr_cry_11 : std_logic;
signal \ctrZ0Z_13\ : std_logic;
signal ctr_cry_12 : std_logic;
signal \ctrZ0Z_14\ : std_logic;
signal ctr_cry_13 : std_logic;
signal \ctrZ0Z_15\ : std_logic;
signal ctr_cry_14 : std_logic;
signal ctr_cry_15 : std_logic;
signal \ctrZ0Z_16\ : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal \ctrZ0Z_17\ : std_logic;
signal ctr_cry_16 : std_logic;
signal ctr_cry_17 : std_logic;
signal \ctrZ0Z_18\ : std_logic;
signal \N_412_i\ : std_logic;
signal \p_vLED_cl_iZ0Z_0\ : std_logic;
signal \N_429_i\ : std_logic;
signal \p_vLED_cl_6_iZ0Z_0\ : std_logic;
signal \N_425_i\ : std_logic;
signal \p_vLED_cl_8_iZ0Z_0\ : std_logic;
signal \N_424_i\ : std_logic;
signal \p_vLED_cl_3_iZ0Z_0\ : std_logic;
signal \N_422_i\ : std_logic;
signal \N_58_cascade_\ : std_logic;
signal \p_vLED_cl_1_iZ0Z_0\ : std_logic;
signal \N_423_i\ : std_logic;
signal \ballXZ0Z_1\ : std_logic;
signal \ballXZ0Z_2\ : std_logic;
signal \ballXZ0Z_0\ : std_logic;
signal \p_hLED52_NE_0\ : std_logic;
signal \N_70_i\ : std_logic;
signal \ballXZ0Z_3\ : std_logic;
signal \N_410_i\ : std_logic;
signal \p_hLED_cl_6_iZ0Z_0\ : std_logic;
signal \p_vLED_cl_4_iZ0Z_0\ : std_logic;
signal \N_427_i\ : std_logic;
signal \p_vLED_cl_7_iZ0Z_0\ : std_logic;
signal \N_426_i\ : std_logic;
signal \N_414_i\ : std_logic;
signal \p_vLED_cl_5_iZ0Z_0\ : std_logic;
signal \N_421_i\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \p_hLED_cl_7_iZ0Z_0\ : std_logic;
signal \p_hLED_cl_iZ0Z_0\ : std_logic;
signal \N_58\ : std_logic;
signal \p_hLED_cl_14_iZ0Z_0\ : std_logic;
signal \N_406_i\ : std_logic;
signal \p_hLED_cl_4_iZ0Z_0\ : std_logic;
signal \N_408_i\ : std_logic;
signal \N_407_i\ : std_logic;
signal \p_hLED_cl_2_iZ0Z_0\ : std_logic;
signal \N_409_i\ : std_logic;
signal \p_hLED_cl_3_iZ0Z_0\ : std_logic;
signal \hIndexZ0Z_3\ : std_logic;
signal \hIndexZ0Z_2\ : std_logic;
signal \hIndexZ0Z_1\ : std_logic;
signal \hIndexZ0Z_0\ : std_logic;
signal p_clk12_c_g : std_logic;
signal \p_hLED52\ : std_logic;
signal \p_hLED_cl_13_iZ0Z_0\ : std_logic;
signal \N_416_i\ : std_logic;
signal \p_hLED_cl_8_iZ0Z_0\ : std_logic;
signal \N_411_i\ : std_logic;
signal \p_hLED_cl_10_iZ0Z_0\ : std_logic;
signal \N_417_i\ : std_logic;
signal \p_hLED_cl_9_iZ0Z_0\ : std_logic;
signal \N_418_i\ : std_logic;
signal \p_hLED_cl_1_iZ0Z_0\ : std_logic;
signal \N_413_i\ : std_logic;
signal \p_hLED_cl_11_iZ0Z_0\ : std_logic;
signal \N_420_i\ : std_logic;
signal \p_hLED_cl_12_iZ0Z_0\ : std_logic;
signal \N_415_i\ : std_logic;
signal \p_hLED_cl_5_iZ0Z_0\ : std_logic;
signal \N_419_i\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal p_clk12_wire : std_logic;
signal \p_vLED_wire\ : std_logic_vector(9 downto 0);
signal \p_hLED_wire\ : std_logic_vector(14 downto 0);

begin
    p_clk12_wire <= p_clk12;
    p_vLED <= \p_vLED_wire\;
    p_hLED <= \p_hLED_wire\;

    \p_clk12_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__3965\,
            GLOBALBUFFEROUTPUT => p_clk12_c_g
        );

    \p_clk12_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__3967\,
            DIN => \N__3966\,
            DOUT => \N__3965\,
            PACKAGEPIN => p_clk12_wire
        );

    \p_clk12_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3967\,
            PADOUT => \N__3966\,
            PADIN => \N__3965\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \p_vLED_obuft_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__3956\,
            DIN => \N__3955\,
            DOUT => \N__3954\,
            PACKAGEPIN => \p_vLED_wire\(0)
        );

    \p_vLED_obuft_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3956\,
            PADOUT => \N__3955\,
            PADIN => \N__3954\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2851\,
            DIN0 => OPEN,
            DOUT0 => \N__3063\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \p_hLED_obuft_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__3947\,
            DIN => \N__3946\,
            DOUT => \N__3945\,
            PACKAGEPIN => \p_hLED_wire\(2)
        );

    \p_hLED_obuft_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3947\,
            PADOUT => \N__3946\,
            PADIN => \N__3945\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2941\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \p_hLED_obuft_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__3938\,
            DIN => \N__3937\,
            DOUT => \N__3936\,
            PACKAGEPIN => \p_hLED_wire\(5)
        );

    \p_hLED_obuft_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3938\,
            PADOUT => \N__3937\,
            PADIN => \N__3936\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3079\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \p_hLED_obuft_10_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__3929\,
            DIN => \N__3928\,
            DOUT => \N__3927\,
            PACKAGEPIN => \p_hLED_wire\(10)
        );

    \p_hLED_obuft_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3929\,
            PADOUT => \N__3928\,
            PADIN => \N__3927\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3097\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \p_vLED_obuft_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__3920\,
            DIN => \N__3919\,
            DOUT => \N__3918\,
            PACKAGEPIN => \p_vLED_wire\(7)
        );

    \p_vLED_obuft_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3920\,
            PADOUT => \N__3919\,
            PADIN => \N__3918\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__1873\,
            DIN0 => OPEN,
            DOUT0 => \N__3072\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \p_vLED_obuft_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__3911\,
            DIN => \N__3910\,
            DOUT => \N__3909\,
            PACKAGEPIN => \p_vLED_wire\(2)
        );

    \p_vLED_obuft_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3911\,
            PADOUT => \N__3910\,
            PADIN => \N__3909\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2821\,
            DIN0 => OPEN,
            DOUT0 => \N__3030\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \p_vLED_obuft_9_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__3902\,
            DIN => \N__3901\,
            DOUT => \N__3900\,
            PACKAGEPIN => \p_vLED_wire\(9)
        );

    \p_vLED_obuft_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3902\,
            PADOUT => \N__3901\,
            PADIN => \N__3900\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__1882\,
            DIN0 => OPEN,
            DOUT0 => \N__3070\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \p_hLED_obuft_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__3893\,
            DIN => \N__3892\,
            DOUT => \N__3891\,
            PACKAGEPIN => \p_hLED_wire\(0)
        );

    \p_hLED_obuft_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3893\,
            PADOUT => \N__3892\,
            PADIN => \N__3891\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2953\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \p_vLED_obuft_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__3884\,
            DIN => \N__3883\,
            DOUT => \N__3882\,
            PACKAGEPIN => \p_vLED_wire\(1)
        );

    \p_vLED_obuft_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3884\,
            PADOUT => \N__3883\,
            PADIN => \N__3882\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2551\,
            DIN0 => OPEN,
            DOUT0 => \N__3031\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \p_hLED_obuft_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__3875\,
            DIN => \N__3874\,
            DOUT => \N__3873\,
            PACKAGEPIN => \p_hLED_wire\(7)
        );

    \p_hLED_obuft_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3875\,
            PADOUT => \N__3874\,
            PADIN => \N__3873\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3664\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \p_hLED_obuft_12_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__3866\,
            DIN => \N__3865\,
            DOUT => \N__3864\,
            PACKAGEPIN => \p_hLED_wire\(12)
        );

    \p_hLED_obuft_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3866\,
            PADOUT => \N__3865\,
            PADIN => \N__3864\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3691\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \p_hLED_obuft_8_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__3857\,
            DIN => \N__3856\,
            DOUT => \N__3855\,
            PACKAGEPIN => \p_hLED_wire\(8)
        );

    \p_hLED_obuft_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3857\,
            PADOUT => \N__3856\,
            PADIN => \N__3855\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2872\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \p_vLED_obuft_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__3848\,
            DIN => \N__3847\,
            DOUT => \N__3846\,
            PACKAGEPIN => \p_vLED_wire\(5)
        );

    \p_vLED_obuft_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3848\,
            PADOUT => \N__3847\,
            PADIN => \N__3846\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2878\,
            DIN0 => OPEN,
            DOUT0 => \N__3062\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \p_hLED_obuft_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__3839\,
            DIN => \N__3838\,
            DOUT => \N__3837\,
            PACKAGEPIN => \p_hLED_wire\(3)
        );

    \p_hLED_obuft_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3839\,
            PADOUT => \N__3838\,
            PADIN => \N__3837\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3598\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \p_hLED_obuft_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__3830\,
            DIN => \N__3829\,
            DOUT => \N__3828\,
            PACKAGEPIN => \p_hLED_wire\(6)
        );

    \p_hLED_obuft_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3830\,
            PADOUT => \N__3829\,
            PADIN => \N__3828\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2632\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \p_hLED_obuft_13_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__3821\,
            DIN => \N__3820\,
            DOUT => \N__3819\,
            PACKAGEPIN => \p_hLED_wire\(13)
        );

    \p_hLED_obuft_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3821\,
            PADOUT => \N__3820\,
            PADIN => \N__3819\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3610\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \p_vLED_obuft_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__3812\,
            DIN => \N__3811\,
            DOUT => \N__3810\,
            PACKAGEPIN => \p_vLED_wire\(4)
        );

    \p_vLED_obuft_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3812\,
            PADOUT => \N__3811\,
            PADIN => \N__3810\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2587\,
            DIN0 => OPEN,
            DOUT0 => \N__3028\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \p_vLED_obuft_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__3803\,
            DIN => \N__3802\,
            DOUT => \N__3801\,
            PACKAGEPIN => \p_vLED_wire\(3)
        );

    \p_vLED_obuft_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3803\,
            PADOUT => \N__3802\,
            PADIN => \N__3801\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2569\,
            DIN0 => OPEN,
            DOUT0 => \N__3029\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \p_hLED_obuft_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__3794\,
            DIN => \N__3793\,
            DOUT => \N__3792\,
            PACKAGEPIN => \p_hLED_wire\(1)
        );

    \p_hLED_obuft_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3794\,
            PADOUT => \N__3793\,
            PADIN => \N__3792\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2935\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \p_hLED_obuft_14_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__3785\,
            DIN => \N__3784\,
            DOUT => \N__3783\,
            PACKAGEPIN => \p_hLED_wire\(14)
        );

    \p_hLED_obuft_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3785\,
            PADOUT => \N__3784\,
            PADIN => \N__3783\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3649\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \p_hLED_obuft_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__3776\,
            DIN => \N__3775\,
            DOUT => \N__3774\,
            PACKAGEPIN => \p_hLED_wire\(4)
        );

    \p_hLED_obuft_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3776\,
            PADOUT => \N__3775\,
            PADIN => \N__3774\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2929\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \p_hLED_obuft_11_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__3767\,
            DIN => \N__3766\,
            DOUT => \N__3765\,
            PACKAGEPIN => \p_hLED_wire\(11)
        );

    \p_hLED_obuft_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3767\,
            PADOUT => \N__3766\,
            PADIN => \N__3765\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3715\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \p_vLED_obuft_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__3758\,
            DIN => \N__3757\,
            DOUT => \N__3756\,
            PACKAGEPIN => \p_vLED_wire\(6)
        );

    \p_vLED_obuft_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3758\,
            PADOUT => \N__3757\,
            PADIN => \N__3756\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2896\,
            DIN0 => OPEN,
            DOUT0 => \N__3073\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \p_hLED_obuft_9_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__3749\,
            DIN => \N__3748\,
            DOUT => \N__3747\,
            PACKAGEPIN => \p_hLED_wire\(9)
        );

    \p_hLED_obuft_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3749\,
            PADOUT => \N__3748\,
            PADIN => \N__3747\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3625\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \p_vLED_obuft_8_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__3740\,
            DIN => \N__3739\,
            DOUT => \N__3738\,
            PACKAGEPIN => \p_vLED_wire\(8)
        );

    \p_vLED_obuft_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__3740\,
            PADOUT => \N__3739\,
            PADIN => \N__3738\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2608\,
            DIN0 => OPEN,
            DOUT0 => \N__3071\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__830\ : InMux
    port map (
            O => \N__3721\,
            I => \N__3718\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__3718\,
            I => \p_hLED_cl_10_iZ0Z_0\
        );

    \I__828\ : IoInMux
    port map (
            O => \N__3715\,
            I => \N__3712\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__3712\,
            I => \N__3709\
        );

    \I__826\ : Span4Mux_s1_h
    port map (
            O => \N__3709\,
            I => \N__3706\
        );

    \I__825\ : Span4Mux_v
    port map (
            O => \N__3706\,
            I => \N__3703\
        );

    \I__824\ : Odrv4
    port map (
            O => \N__3703\,
            I => \N_417_i\
        );

    \I__823\ : InMux
    port map (
            O => \N__3700\,
            I => \N__3697\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__3697\,
            I => \N__3694\
        );

    \I__821\ : Odrv12
    port map (
            O => \N__3694\,
            I => \p_hLED_cl_9_iZ0Z_0\
        );

    \I__820\ : IoInMux
    port map (
            O => \N__3691\,
            I => \N__3688\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__3688\,
            I => \N__3685\
        );

    \I__818\ : IoSpan4Mux
    port map (
            O => \N__3685\,
            I => \N__3682\
        );

    \I__817\ : Span4Mux_s3_v
    port map (
            O => \N__3682\,
            I => \N__3679\
        );

    \I__816\ : Odrv4
    port map (
            O => \N__3679\,
            I => \N_418_i\
        );

    \I__815\ : InMux
    port map (
            O => \N__3676\,
            I => \N__3673\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__3673\,
            I => \N__3670\
        );

    \I__813\ : Span12Mux_s9_v
    port map (
            O => \N__3670\,
            I => \N__3667\
        );

    \I__812\ : Odrv12
    port map (
            O => \N__3667\,
            I => \p_hLED_cl_1_iZ0Z_0\
        );

    \I__811\ : IoInMux
    port map (
            O => \N__3664\,
            I => \N__3661\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__3661\,
            I => \N_413_i\
        );

    \I__809\ : InMux
    port map (
            O => \N__3658\,
            I => \N__3655\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__3655\,
            I => \N__3652\
        );

    \I__807\ : Odrv12
    port map (
            O => \N__3652\,
            I => \p_hLED_cl_11_iZ0Z_0\
        );

    \I__806\ : IoInMux
    port map (
            O => \N__3649\,
            I => \N__3646\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__3646\,
            I => \N__3643\
        );

    \I__804\ : Span4Mux_s0_h
    port map (
            O => \N__3643\,
            I => \N__3640\
        );

    \I__803\ : Odrv4
    port map (
            O => \N__3640\,
            I => \N_420_i\
        );

    \I__802\ : InMux
    port map (
            O => \N__3637\,
            I => \N__3634\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__3634\,
            I => \N__3631\
        );

    \I__800\ : Span4Mux_v
    port map (
            O => \N__3631\,
            I => \N__3628\
        );

    \I__799\ : Odrv4
    port map (
            O => \N__3628\,
            I => \p_hLED_cl_12_iZ0Z_0\
        );

    \I__798\ : IoInMux
    port map (
            O => \N__3625\,
            I => \N__3622\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__3622\,
            I => \N_415_i\
        );

    \I__796\ : InMux
    port map (
            O => \N__3619\,
            I => \N__3616\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__3616\,
            I => \N__3613\
        );

    \I__794\ : Odrv12
    port map (
            O => \N__3613\,
            I => \p_hLED_cl_5_iZ0Z_0\
        );

    \I__793\ : IoInMux
    port map (
            O => \N__3610\,
            I => \N__3607\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__3607\,
            I => \N_419_i\
        );

    \I__791\ : InMux
    port map (
            O => \N__3604\,
            I => \N__3601\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__3601\,
            I => \p_hLED_cl_2_iZ0Z_0\
        );

    \I__789\ : IoInMux
    port map (
            O => \N__3598\,
            I => \N__3595\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__3595\,
            I => \N_409_i\
        );

    \I__787\ : InMux
    port map (
            O => \N__3592\,
            I => \N__3589\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__3589\,
            I => \p_hLED_cl_3_iZ0Z_0\
        );

    \I__785\ : CascadeMux
    port map (
            O => \N__3586\,
            I => \N__3577\
        );

    \I__784\ : InMux
    port map (
            O => \N__3585\,
            I => \N__3550\
        );

    \I__783\ : InMux
    port map (
            O => \N__3584\,
            I => \N__3550\
        );

    \I__782\ : InMux
    port map (
            O => \N__3583\,
            I => \N__3550\
        );

    \I__781\ : InMux
    port map (
            O => \N__3582\,
            I => \N__3550\
        );

    \I__780\ : InMux
    port map (
            O => \N__3581\,
            I => \N__3550\
        );

    \I__779\ : InMux
    port map (
            O => \N__3580\,
            I => \N__3550\
        );

    \I__778\ : InMux
    port map (
            O => \N__3577\,
            I => \N__3547\
        );

    \I__777\ : InMux
    port map (
            O => \N__3576\,
            I => \N__3538\
        );

    \I__776\ : InMux
    port map (
            O => \N__3575\,
            I => \N__3538\
        );

    \I__775\ : InMux
    port map (
            O => \N__3574\,
            I => \N__3538\
        );

    \I__774\ : InMux
    port map (
            O => \N__3573\,
            I => \N__3538\
        );

    \I__773\ : InMux
    port map (
            O => \N__3572\,
            I => \N__3535\
        );

    \I__772\ : InMux
    port map (
            O => \N__3571\,
            I => \N__3526\
        );

    \I__771\ : InMux
    port map (
            O => \N__3570\,
            I => \N__3526\
        );

    \I__770\ : InMux
    port map (
            O => \N__3569\,
            I => \N__3526\
        );

    \I__769\ : InMux
    port map (
            O => \N__3568\,
            I => \N__3526\
        );

    \I__768\ : InMux
    port map (
            O => \N__3567\,
            I => \N__3515\
        );

    \I__767\ : InMux
    port map (
            O => \N__3566\,
            I => \N__3515\
        );

    \I__766\ : InMux
    port map (
            O => \N__3565\,
            I => \N__3515\
        );

    \I__765\ : InMux
    port map (
            O => \N__3564\,
            I => \N__3515\
        );

    \I__764\ : InMux
    port map (
            O => \N__3563\,
            I => \N__3515\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__3550\,
            I => \N__3512\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__3547\,
            I => \N__3509\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__3538\,
            I => \N__3504\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__3535\,
            I => \N__3504\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__3526\,
            I => \hIndexZ0Z_3\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__3515\,
            I => \hIndexZ0Z_3\
        );

    \I__757\ : Odrv4
    port map (
            O => \N__3512\,
            I => \hIndexZ0Z_3\
        );

    \I__756\ : Odrv4
    port map (
            O => \N__3509\,
            I => \hIndexZ0Z_3\
        );

    \I__755\ : Odrv4
    port map (
            O => \N__3504\,
            I => \hIndexZ0Z_3\
        );

    \I__754\ : InMux
    port map (
            O => \N__3493\,
            I => \N__3467\
        );

    \I__753\ : InMux
    port map (
            O => \N__3492\,
            I => \N__3467\
        );

    \I__752\ : InMux
    port map (
            O => \N__3491\,
            I => \N__3467\
        );

    \I__751\ : InMux
    port map (
            O => \N__3490\,
            I => \N__3467\
        );

    \I__750\ : InMux
    port map (
            O => \N__3489\,
            I => \N__3467\
        );

    \I__749\ : InMux
    port map (
            O => \N__3488\,
            I => \N__3467\
        );

    \I__748\ : InMux
    port map (
            O => \N__3487\,
            I => \N__3458\
        );

    \I__747\ : InMux
    port map (
            O => \N__3486\,
            I => \N__3458\
        );

    \I__746\ : InMux
    port map (
            O => \N__3485\,
            I => \N__3458\
        );

    \I__745\ : InMux
    port map (
            O => \N__3484\,
            I => \N__3458\
        );

    \I__744\ : InMux
    port map (
            O => \N__3483\,
            I => \N__3452\
        );

    \I__743\ : InMux
    port map (
            O => \N__3482\,
            I => \N__3444\
        );

    \I__742\ : InMux
    port map (
            O => \N__3481\,
            I => \N__3444\
        );

    \I__741\ : InMux
    port map (
            O => \N__3480\,
            I => \N__3444\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__3467\,
            I => \N__3441\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__3458\,
            I => \N__3438\
        );

    \I__738\ : InMux
    port map (
            O => \N__3457\,
            I => \N__3431\
        );

    \I__737\ : InMux
    port map (
            O => \N__3456\,
            I => \N__3431\
        );

    \I__736\ : InMux
    port map (
            O => \N__3455\,
            I => \N__3431\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__3452\,
            I => \N__3428\
        );

    \I__734\ : InMux
    port map (
            O => \N__3451\,
            I => \N__3425\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__3444\,
            I => \hIndexZ0Z_2\
        );

    \I__732\ : Odrv4
    port map (
            O => \N__3441\,
            I => \hIndexZ0Z_2\
        );

    \I__731\ : Odrv4
    port map (
            O => \N__3438\,
            I => \hIndexZ0Z_2\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__3431\,
            I => \hIndexZ0Z_2\
        );

    \I__729\ : Odrv12
    port map (
            O => \N__3428\,
            I => \hIndexZ0Z_2\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__3425\,
            I => \hIndexZ0Z_2\
        );

    \I__727\ : CascadeMux
    port map (
            O => \N__3412\,
            I => \N__3396\
        );

    \I__726\ : CascadeMux
    port map (
            O => \N__3411\,
            I => \N__3393\
        );

    \I__725\ : CascadeMux
    port map (
            O => \N__3410\,
            I => \N__3390\
        );

    \I__724\ : CascadeMux
    port map (
            O => \N__3409\,
            I => \N__3387\
        );

    \I__723\ : CascadeMux
    port map (
            O => \N__3408\,
            I => \N__3384\
        );

    \I__722\ : CascadeMux
    port map (
            O => \N__3407\,
            I => \N__3381\
        );

    \I__721\ : CascadeMux
    port map (
            O => \N__3406\,
            I => \N__3376\
        );

    \I__720\ : CascadeMux
    port map (
            O => \N__3405\,
            I => \N__3373\
        );

    \I__719\ : CascadeMux
    port map (
            O => \N__3404\,
            I => \N__3370\
        );

    \I__718\ : CascadeMux
    port map (
            O => \N__3403\,
            I => \N__3367\
        );

    \I__717\ : CascadeMux
    port map (
            O => \N__3402\,
            I => \N__3364\
        );

    \I__716\ : InMux
    port map (
            O => \N__3401\,
            I => \N__3351\
        );

    \I__715\ : InMux
    port map (
            O => \N__3400\,
            I => \N__3351\
        );

    \I__714\ : InMux
    port map (
            O => \N__3399\,
            I => \N__3351\
        );

    \I__713\ : InMux
    port map (
            O => \N__3396\,
            I => \N__3351\
        );

    \I__712\ : InMux
    port map (
            O => \N__3393\,
            I => \N__3351\
        );

    \I__711\ : InMux
    port map (
            O => \N__3390\,
            I => \N__3351\
        );

    \I__710\ : InMux
    port map (
            O => \N__3387\,
            I => \N__3342\
        );

    \I__709\ : InMux
    port map (
            O => \N__3384\,
            I => \N__3342\
        );

    \I__708\ : InMux
    port map (
            O => \N__3381\,
            I => \N__3342\
        );

    \I__707\ : InMux
    port map (
            O => \N__3380\,
            I => \N__3342\
        );

    \I__706\ : InMux
    port map (
            O => \N__3379\,
            I => \N__3338\
        );

    \I__705\ : InMux
    port map (
            O => \N__3376\,
            I => \N__3334\
        );

    \I__704\ : InMux
    port map (
            O => \N__3373\,
            I => \N__3329\
        );

    \I__703\ : InMux
    port map (
            O => \N__3370\,
            I => \N__3329\
        );

    \I__702\ : InMux
    port map (
            O => \N__3367\,
            I => \N__3324\
        );

    \I__701\ : InMux
    port map (
            O => \N__3364\,
            I => \N__3324\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__3351\,
            I => \N__3321\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__3342\,
            I => \N__3318\
        );

    \I__698\ : InMux
    port map (
            O => \N__3341\,
            I => \N__3315\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__3338\,
            I => \N__3312\
        );

    \I__696\ : InMux
    port map (
            O => \N__3337\,
            I => \N__3309\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__3334\,
            I => \hIndexZ0Z_1\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__3329\,
            I => \hIndexZ0Z_1\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__3324\,
            I => \hIndexZ0Z_1\
        );

    \I__692\ : Odrv4
    port map (
            O => \N__3321\,
            I => \hIndexZ0Z_1\
        );

    \I__691\ : Odrv4
    port map (
            O => \N__3318\,
            I => \hIndexZ0Z_1\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__3315\,
            I => \hIndexZ0Z_1\
        );

    \I__689\ : Odrv4
    port map (
            O => \N__3312\,
            I => \hIndexZ0Z_1\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__3309\,
            I => \hIndexZ0Z_1\
        );

    \I__687\ : CascadeMux
    port map (
            O => \N__3292\,
            I => \N__3286\
        );

    \I__686\ : CascadeMux
    port map (
            O => \N__3291\,
            I => \N__3277\
        );

    \I__685\ : CascadeMux
    port map (
            O => \N__3290\,
            I => \N__3274\
        );

    \I__684\ : CascadeMux
    port map (
            O => \N__3289\,
            I => \N__3271\
        );

    \I__683\ : InMux
    port map (
            O => \N__3286\,
            I => \N__3262\
        );

    \I__682\ : InMux
    port map (
            O => \N__3285\,
            I => \N__3262\
        );

    \I__681\ : InMux
    port map (
            O => \N__3284\,
            I => \N__3262\
        );

    \I__680\ : InMux
    port map (
            O => \N__3283\,
            I => \N__3262\
        );

    \I__679\ : InMux
    port map (
            O => \N__3282\,
            I => \N__3249\
        );

    \I__678\ : InMux
    port map (
            O => \N__3281\,
            I => \N__3249\
        );

    \I__677\ : InMux
    port map (
            O => \N__3280\,
            I => \N__3249\
        );

    \I__676\ : InMux
    port map (
            O => \N__3277\,
            I => \N__3249\
        );

    \I__675\ : InMux
    port map (
            O => \N__3274\,
            I => \N__3249\
        );

    \I__674\ : InMux
    port map (
            O => \N__3271\,
            I => \N__3249\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__3262\,
            I => \N__3234\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__3249\,
            I => \N__3234\
        );

    \I__671\ : InMux
    port map (
            O => \N__3248\,
            I => \N__3231\
        );

    \I__670\ : InMux
    port map (
            O => \N__3247\,
            I => \N__3225\
        );

    \I__669\ : InMux
    port map (
            O => \N__3246\,
            I => \N__3225\
        );

    \I__668\ : InMux
    port map (
            O => \N__3245\,
            I => \N__3220\
        );

    \I__667\ : InMux
    port map (
            O => \N__3244\,
            I => \N__3220\
        );

    \I__666\ : InMux
    port map (
            O => \N__3243\,
            I => \N__3213\
        );

    \I__665\ : InMux
    port map (
            O => \N__3242\,
            I => \N__3213\
        );

    \I__664\ : InMux
    port map (
            O => \N__3241\,
            I => \N__3213\
        );

    \I__663\ : InMux
    port map (
            O => \N__3240\,
            I => \N__3210\
        );

    \I__662\ : InMux
    port map (
            O => \N__3239\,
            I => \N__3207\
        );

    \I__661\ : Span4Mux_v
    port map (
            O => \N__3234\,
            I => \N__3204\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__3231\,
            I => \N__3201\
        );

    \I__659\ : InMux
    port map (
            O => \N__3230\,
            I => \N__3198\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__3225\,
            I => \hIndexZ0Z_0\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__3220\,
            I => \hIndexZ0Z_0\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__3213\,
            I => \hIndexZ0Z_0\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__3210\,
            I => \hIndexZ0Z_0\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__3207\,
            I => \hIndexZ0Z_0\
        );

    \I__653\ : Odrv4
    port map (
            O => \N__3204\,
            I => \hIndexZ0Z_0\
        );

    \I__652\ : Odrv4
    port map (
            O => \N__3201\,
            I => \hIndexZ0Z_0\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__3198\,
            I => \hIndexZ0Z_0\
        );

    \I__650\ : ClkMux
    port map (
            O => \N__3181\,
            I => \N__3142\
        );

    \I__649\ : ClkMux
    port map (
            O => \N__3180\,
            I => \N__3142\
        );

    \I__648\ : ClkMux
    port map (
            O => \N__3179\,
            I => \N__3142\
        );

    \I__647\ : ClkMux
    port map (
            O => \N__3178\,
            I => \N__3142\
        );

    \I__646\ : ClkMux
    port map (
            O => \N__3177\,
            I => \N__3142\
        );

    \I__645\ : ClkMux
    port map (
            O => \N__3176\,
            I => \N__3142\
        );

    \I__644\ : ClkMux
    port map (
            O => \N__3175\,
            I => \N__3142\
        );

    \I__643\ : ClkMux
    port map (
            O => \N__3174\,
            I => \N__3142\
        );

    \I__642\ : ClkMux
    port map (
            O => \N__3173\,
            I => \N__3142\
        );

    \I__641\ : ClkMux
    port map (
            O => \N__3172\,
            I => \N__3142\
        );

    \I__640\ : ClkMux
    port map (
            O => \N__3171\,
            I => \N__3142\
        );

    \I__639\ : ClkMux
    port map (
            O => \N__3170\,
            I => \N__3142\
        );

    \I__638\ : ClkMux
    port map (
            O => \N__3169\,
            I => \N__3142\
        );

    \I__637\ : GlobalMux
    port map (
            O => \N__3142\,
            I => \N__3139\
        );

    \I__636\ : gio2CtrlBuf
    port map (
            O => \N__3139\,
            I => p_clk12_c_g
        );

    \I__635\ : CEMux
    port map (
            O => \N__3136\,
            I => \N__3132\
        );

    \I__634\ : CEMux
    port map (
            O => \N__3135\,
            I => \N__3128\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__3132\,
            I => \N__3125\
        );

    \I__632\ : CEMux
    port map (
            O => \N__3131\,
            I => \N__3122\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__3128\,
            I => \N__3119\
        );

    \I__630\ : Span4Mux_v
    port map (
            O => \N__3125\,
            I => \N__3114\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__3122\,
            I => \N__3114\
        );

    \I__628\ : Span4Mux_v
    port map (
            O => \N__3119\,
            I => \N__3109\
        );

    \I__627\ : Span4Mux_s0_h
    port map (
            O => \N__3114\,
            I => \N__3109\
        );

    \I__626\ : Span4Mux_h
    port map (
            O => \N__3109\,
            I => \N__3106\
        );

    \I__625\ : Odrv4
    port map (
            O => \N__3106\,
            I => \p_hLED52\
        );

    \I__624\ : InMux
    port map (
            O => \N__3103\,
            I => \N__3100\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__3100\,
            I => \p_hLED_cl_13_iZ0Z_0\
        );

    \I__622\ : IoInMux
    port map (
            O => \N__3097\,
            I => \N__3094\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__3094\,
            I => \N__3091\
        );

    \I__620\ : Span4Mux_s0_h
    port map (
            O => \N__3091\,
            I => \N__3088\
        );

    \I__619\ : Odrv4
    port map (
            O => \N__3088\,
            I => \N_416_i\
        );

    \I__618\ : InMux
    port map (
            O => \N__3085\,
            I => \N__3082\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__3082\,
            I => \p_hLED_cl_8_iZ0Z_0\
        );

    \I__616\ : IoInMux
    port map (
            O => \N__3079\,
            I => \N__3076\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__3076\,
            I => \N_411_i\
        );

    \I__614\ : IoInMux
    port map (
            O => \N__3073\,
            I => \N__3067\
        );

    \I__613\ : IoInMux
    port map (
            O => \N__3072\,
            I => \N__3064\
        );

    \I__612\ : IoInMux
    port map (
            O => \N__3071\,
            I => \N__3059\
        );

    \I__611\ : IoInMux
    port map (
            O => \N__3070\,
            I => \N__3056\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__3067\,
            I => \N__3051\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__3064\,
            I => \N__3051\
        );

    \I__608\ : IoInMux
    port map (
            O => \N__3063\,
            I => \N__3048\
        );

    \I__607\ : IoInMux
    port map (
            O => \N__3062\,
            I => \N__3045\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__3059\,
            I => \N__3038\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__3056\,
            I => \N__3038\
        );

    \I__604\ : IoSpan4Mux
    port map (
            O => \N__3051\,
            I => \N__3038\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__3048\,
            I => \N__3035\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__3045\,
            I => \N__3032\
        );

    \I__601\ : Span4Mux_s0_h
    port map (
            O => \N__3038\,
            I => \N__3025\
        );

    \I__600\ : Span4Mux_s0_h
    port map (
            O => \N__3035\,
            I => \N__3020\
        );

    \I__599\ : Span4Mux_s0_h
    port map (
            O => \N__3032\,
            I => \N__3020\
        );

    \I__598\ : IoInMux
    port map (
            O => \N__3031\,
            I => \N__3017\
        );

    \I__597\ : IoInMux
    port map (
            O => \N__3030\,
            I => \N__3014\
        );

    \I__596\ : IoInMux
    port map (
            O => \N__3029\,
            I => \N__3011\
        );

    \I__595\ : IoInMux
    port map (
            O => \N__3028\,
            I => \N__3008\
        );

    \I__594\ : Odrv4
    port map (
            O => \N__3025\,
            I => \CONSTANT_ONE_NET\
        );

    \I__593\ : Odrv4
    port map (
            O => \N__3020\,
            I => \CONSTANT_ONE_NET\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__3017\,
            I => \CONSTANT_ONE_NET\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__3014\,
            I => \CONSTANT_ONE_NET\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__3011\,
            I => \CONSTANT_ONE_NET\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__3008\,
            I => \CONSTANT_ONE_NET\
        );

    \I__588\ : InMux
    port map (
            O => \N__2995\,
            I => \N__2992\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__2992\,
            I => \N__2989\
        );

    \I__586\ : Span4Mux_v
    port map (
            O => \N__2989\,
            I => \N__2986\
        );

    \I__585\ : Odrv4
    port map (
            O => \N__2986\,
            I => \p_hLED_cl_7_iZ0Z_0\
        );

    \I__584\ : InMux
    port map (
            O => \N__2983\,
            I => \N__2980\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__2980\,
            I => \N__2977\
        );

    \I__582\ : Odrv4
    port map (
            O => \N__2977\,
            I => \p_hLED_cl_iZ0Z_0\
        );

    \I__581\ : InMux
    port map (
            O => \N__2974\,
            I => \N__2967\
        );

    \I__580\ : InMux
    port map (
            O => \N__2973\,
            I => \N__2967\
        );

    \I__579\ : InMux
    port map (
            O => \N__2972\,
            I => \N__2964\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__2967\,
            I => \N_58\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__2964\,
            I => \N_58\
        );

    \I__576\ : InMux
    port map (
            O => \N__2959\,
            I => \N__2956\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__2956\,
            I => \p_hLED_cl_14_iZ0Z_0\
        );

    \I__574\ : IoInMux
    port map (
            O => \N__2953\,
            I => \N__2950\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__2950\,
            I => \N_406_i\
        );

    \I__572\ : InMux
    port map (
            O => \N__2947\,
            I => \N__2944\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__2944\,
            I => \p_hLED_cl_4_iZ0Z_0\
        );

    \I__570\ : IoInMux
    port map (
            O => \N__2941\,
            I => \N__2938\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__2938\,
            I => \N_408_i\
        );

    \I__568\ : IoInMux
    port map (
            O => \N__2935\,
            I => \N__2932\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__2932\,
            I => \N_407_i\
        );

    \I__566\ : IoInMux
    port map (
            O => \N__2929\,
            I => \N__2926\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__2926\,
            I => \N__2923\
        );

    \I__564\ : IoSpan4Mux
    port map (
            O => \N__2923\,
            I => \N__2920\
        );

    \I__563\ : Span4Mux_s1_h
    port map (
            O => \N__2920\,
            I => \N__2917\
        );

    \I__562\ : Odrv4
    port map (
            O => \N__2917\,
            I => \N_410_i\
        );

    \I__561\ : InMux
    port map (
            O => \N__2914\,
            I => \N__2911\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__2911\,
            I => \p_hLED_cl_6_iZ0Z_0\
        );

    \I__559\ : InMux
    port map (
            O => \N__2908\,
            I => \N__2905\
        );

    \I__558\ : LocalMux
    port map (
            O => \N__2905\,
            I => \N__2902\
        );

    \I__557\ : Span4Mux_s3_v
    port map (
            O => \N__2902\,
            I => \N__2899\
        );

    \I__556\ : Odrv4
    port map (
            O => \N__2899\,
            I => \p_vLED_cl_4_iZ0Z_0\
        );

    \I__555\ : IoInMux
    port map (
            O => \N__2896\,
            I => \N__2893\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__2893\,
            I => \N_427_i\
        );

    \I__553\ : InMux
    port map (
            O => \N__2890\,
            I => \N__2887\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__2887\,
            I => \N__2884\
        );

    \I__551\ : Span4Mux_s3_h
    port map (
            O => \N__2884\,
            I => \N__2881\
        );

    \I__550\ : Odrv4
    port map (
            O => \N__2881\,
            I => \p_vLED_cl_7_iZ0Z_0\
        );

    \I__549\ : IoInMux
    port map (
            O => \N__2878\,
            I => \N__2875\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__2875\,
            I => \N_426_i\
        );

    \I__547\ : IoInMux
    port map (
            O => \N__2872\,
            I => \N__2869\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__2869\,
            I => \N__2866\
        );

    \I__545\ : Span4Mux_s3_v
    port map (
            O => \N__2866\,
            I => \N__2863\
        );

    \I__544\ : Odrv4
    port map (
            O => \N__2863\,
            I => \N_414_i\
        );

    \I__543\ : InMux
    port map (
            O => \N__2860\,
            I => \N__2857\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__2857\,
            I => \N__2854\
        );

    \I__541\ : Odrv12
    port map (
            O => \N__2854\,
            I => \p_vLED_cl_5_iZ0Z_0\
        );

    \I__540\ : IoInMux
    port map (
            O => \N__2851\,
            I => \N__2848\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__2848\,
            I => \N__2845\
        );

    \I__538\ : Span4Mux_s0_h
    port map (
            O => \N__2845\,
            I => \N__2842\
        );

    \I__537\ : Sp12to4
    port map (
            O => \N__2842\,
            I => \N__2839\
        );

    \I__536\ : Odrv12
    port map (
            O => \N__2839\,
            I => \N_421_i\
        );

    \I__535\ : CascadeMux
    port map (
            O => \N__2836\,
            I => \N_58_cascade_\
        );

    \I__534\ : InMux
    port map (
            O => \N__2833\,
            I => \N__2830\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__2830\,
            I => \N__2827\
        );

    \I__532\ : Span4Mux_v
    port map (
            O => \N__2827\,
            I => \N__2824\
        );

    \I__531\ : Odrv4
    port map (
            O => \N__2824\,
            I => \p_vLED_cl_1_iZ0Z_0\
        );

    \I__530\ : IoInMux
    port map (
            O => \N__2821\,
            I => \N__2818\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__2818\,
            I => \N__2815\
        );

    \I__528\ : Odrv12
    port map (
            O => \N__2815\,
            I => \N_423_i\
        );

    \I__527\ : InMux
    port map (
            O => \N__2812\,
            I => \N__2807\
        );

    \I__526\ : InMux
    port map (
            O => \N__2811\,
            I => \N__2804\
        );

    \I__525\ : InMux
    port map (
            O => \N__2810\,
            I => \N__2801\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__2807\,
            I => \N__2798\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__2804\,
            I => \ballXZ0Z_1\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__2801\,
            I => \ballXZ0Z_1\
        );

    \I__521\ : Odrv12
    port map (
            O => \N__2798\,
            I => \ballXZ0Z_1\
        );

    \I__520\ : CascadeMux
    port map (
            O => \N__2791\,
            I => \N__2787\
        );

    \I__519\ : CascadeMux
    port map (
            O => \N__2790\,
            I => \N__2783\
        );

    \I__518\ : InMux
    port map (
            O => \N__2787\,
            I => \N__2780\
        );

    \I__517\ : InMux
    port map (
            O => \N__2786\,
            I => \N__2777\
        );

    \I__516\ : InMux
    port map (
            O => \N__2783\,
            I => \N__2774\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__2780\,
            I => \N__2771\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__2777\,
            I => \ballXZ0Z_2\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__2774\,
            I => \ballXZ0Z_2\
        );

    \I__512\ : Odrv12
    port map (
            O => \N__2771\,
            I => \ballXZ0Z_2\
        );

    \I__511\ : InMux
    port map (
            O => \N__2764\,
            I => \N__2759\
        );

    \I__510\ : InMux
    port map (
            O => \N__2763\,
            I => \N__2754\
        );

    \I__509\ : InMux
    port map (
            O => \N__2762\,
            I => \N__2754\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__2759\,
            I => \N__2751\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__2754\,
            I => \ballXZ0Z_0\
        );

    \I__506\ : Odrv12
    port map (
            O => \N__2751\,
            I => \ballXZ0Z_0\
        );

    \I__505\ : InMux
    port map (
            O => \N__2746\,
            I => \N__2743\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__2743\,
            I => \p_hLED52_NE_0\
        );

    \I__503\ : InMux
    port map (
            O => \N__2740\,
            I => \N__2737\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__2737\,
            I => \N_70_i\
        );

    \I__501\ : CascadeMux
    port map (
            O => \N__2734\,
            I => \N__2731\
        );

    \I__500\ : InMux
    port map (
            O => \N__2731\,
            I => \N__2728\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__2728\,
            I => \N__2723\
        );

    \I__498\ : InMux
    port map (
            O => \N__2727\,
            I => \N__2718\
        );

    \I__497\ : InMux
    port map (
            O => \N__2726\,
            I => \N__2718\
        );

    \I__496\ : Span4Mux_h
    port map (
            O => \N__2723\,
            I => \N__2715\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__2718\,
            I => \ballXZ0Z_3\
        );

    \I__494\ : Odrv4
    port map (
            O => \N__2715\,
            I => \ballXZ0Z_3\
        );

    \I__493\ : InMux
    port map (
            O => \N__2710\,
            I => \N__2706\
        );

    \I__492\ : InMux
    port map (
            O => \N__2709\,
            I => \N__2703\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__2706\,
            I => \N__2700\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__2703\,
            I => \ctrZ0Z_15\
        );

    \I__489\ : Odrv4
    port map (
            O => \N__2700\,
            I => \ctrZ0Z_15\
        );

    \I__488\ : InMux
    port map (
            O => \N__2695\,
            I => ctr_cry_14
        );

    \I__487\ : InMux
    port map (
            O => \N__2692\,
            I => \N__2689\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__2689\,
            I => \N__2685\
        );

    \I__485\ : InMux
    port map (
            O => \N__2688\,
            I => \N__2682\
        );

    \I__484\ : Span4Mux_h
    port map (
            O => \N__2685\,
            I => \N__2679\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__2682\,
            I => \ctrZ0Z_16\
        );

    \I__482\ : Odrv4
    port map (
            O => \N__2679\,
            I => \ctrZ0Z_16\
        );

    \I__481\ : InMux
    port map (
            O => \N__2674\,
            I => \bfn_9_9_0_\
        );

    \I__480\ : InMux
    port map (
            O => \N__2671\,
            I => \N__2668\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__2668\,
            I => \N__2664\
        );

    \I__478\ : InMux
    port map (
            O => \N__2667\,
            I => \N__2661\
        );

    \I__477\ : Span4Mux_h
    port map (
            O => \N__2664\,
            I => \N__2658\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__2661\,
            I => \ctrZ0Z_17\
        );

    \I__475\ : Odrv4
    port map (
            O => \N__2658\,
            I => \ctrZ0Z_17\
        );

    \I__474\ : InMux
    port map (
            O => \N__2653\,
            I => ctr_cry_16
        );

    \I__473\ : InMux
    port map (
            O => \N__2650\,
            I => ctr_cry_17
        );

    \I__472\ : InMux
    port map (
            O => \N__2647\,
            I => \N__2643\
        );

    \I__471\ : InMux
    port map (
            O => \N__2646\,
            I => \N__2640\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__2643\,
            I => \N__2637\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__2640\,
            I => \ctrZ0Z_18\
        );

    \I__468\ : Odrv4
    port map (
            O => \N__2637\,
            I => \ctrZ0Z_18\
        );

    \I__467\ : IoInMux
    port map (
            O => \N__2632\,
            I => \N__2629\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__2629\,
            I => \N__2626\
        );

    \I__465\ : Span4Mux_s1_v
    port map (
            O => \N__2626\,
            I => \N__2623\
        );

    \I__464\ : Odrv4
    port map (
            O => \N__2623\,
            I => \N_412_i\
        );

    \I__463\ : InMux
    port map (
            O => \N__2620\,
            I => \N__2617\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__2617\,
            I => \N__2614\
        );

    \I__461\ : Span4Mux_s3_v
    port map (
            O => \N__2614\,
            I => \N__2611\
        );

    \I__460\ : Odrv4
    port map (
            O => \N__2611\,
            I => \p_vLED_cl_iZ0Z_0\
        );

    \I__459\ : IoInMux
    port map (
            O => \N__2608\,
            I => \N__2605\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__2605\,
            I => \N__2602\
        );

    \I__457\ : Span4Mux_s1_h
    port map (
            O => \N__2602\,
            I => \N__2599\
        );

    \I__456\ : Odrv4
    port map (
            O => \N__2599\,
            I => \N_429_i\
        );

    \I__455\ : InMux
    port map (
            O => \N__2596\,
            I => \N__2593\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__2593\,
            I => \N__2590\
        );

    \I__453\ : Odrv4
    port map (
            O => \N__2590\,
            I => \p_vLED_cl_6_iZ0Z_0\
        );

    \I__452\ : IoInMux
    port map (
            O => \N__2587\,
            I => \N__2584\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__2584\,
            I => \N__2581\
        );

    \I__450\ : Odrv4
    port map (
            O => \N__2581\,
            I => \N_425_i\
        );

    \I__449\ : InMux
    port map (
            O => \N__2578\,
            I => \N__2575\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__2575\,
            I => \N__2572\
        );

    \I__447\ : Odrv4
    port map (
            O => \N__2572\,
            I => \p_vLED_cl_8_iZ0Z_0\
        );

    \I__446\ : IoInMux
    port map (
            O => \N__2569\,
            I => \N__2566\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__2566\,
            I => \N__2563\
        );

    \I__444\ : Odrv12
    port map (
            O => \N__2563\,
            I => \N_424_i\
        );

    \I__443\ : InMux
    port map (
            O => \N__2560\,
            I => \N__2557\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__2557\,
            I => \N__2554\
        );

    \I__441\ : Odrv4
    port map (
            O => \N__2554\,
            I => \p_vLED_cl_3_iZ0Z_0\
        );

    \I__440\ : IoInMux
    port map (
            O => \N__2551\,
            I => \N__2548\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__2548\,
            I => \N__2545\
        );

    \I__438\ : IoSpan4Mux
    port map (
            O => \N__2545\,
            I => \N__2542\
        );

    \I__437\ : Odrv4
    port map (
            O => \N__2542\,
            I => \N_422_i\
        );

    \I__436\ : CascadeMux
    port map (
            O => \N__2539\,
            I => \N__2535\
        );

    \I__435\ : InMux
    port map (
            O => \N__2538\,
            I => \N__2532\
        );

    \I__434\ : InMux
    port map (
            O => \N__2535\,
            I => \N__2529\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__2532\,
            I => \N__2524\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__2529\,
            I => \N__2524\
        );

    \I__431\ : Odrv4
    port map (
            O => \N__2524\,
            I => \ctrZ0Z_7\
        );

    \I__430\ : InMux
    port map (
            O => \N__2521\,
            I => ctr_cry_6
        );

    \I__429\ : InMux
    port map (
            O => \N__2518\,
            I => \N__2514\
        );

    \I__428\ : InMux
    port map (
            O => \N__2517\,
            I => \N__2511\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__2514\,
            I => \ctrZ0Z_8\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__2511\,
            I => \ctrZ0Z_8\
        );

    \I__425\ : InMux
    port map (
            O => \N__2506\,
            I => \bfn_9_8_0_\
        );

    \I__424\ : InMux
    port map (
            O => \N__2503\,
            I => \N__2499\
        );

    \I__423\ : InMux
    port map (
            O => \N__2502\,
            I => \N__2496\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__2499\,
            I => \N__2493\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__2496\,
            I => \ctrZ0Z_9\
        );

    \I__420\ : Odrv4
    port map (
            O => \N__2493\,
            I => \ctrZ0Z_9\
        );

    \I__419\ : InMux
    port map (
            O => \N__2488\,
            I => ctr_cry_8
        );

    \I__418\ : InMux
    port map (
            O => \N__2485\,
            I => \N__2481\
        );

    \I__417\ : InMux
    port map (
            O => \N__2484\,
            I => \N__2478\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__2481\,
            I => \ctrZ0Z_10\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__2478\,
            I => \ctrZ0Z_10\
        );

    \I__414\ : InMux
    port map (
            O => \N__2473\,
            I => ctr_cry_9
        );

    \I__413\ : InMux
    port map (
            O => \N__2470\,
            I => \N__2466\
        );

    \I__412\ : InMux
    port map (
            O => \N__2469\,
            I => \N__2463\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__2466\,
            I => \ctrZ0Z_11\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__2463\,
            I => \ctrZ0Z_11\
        );

    \I__409\ : InMux
    port map (
            O => \N__2458\,
            I => ctr_cry_10
        );

    \I__408\ : InMux
    port map (
            O => \N__2455\,
            I => \N__2451\
        );

    \I__407\ : InMux
    port map (
            O => \N__2454\,
            I => \N__2448\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__2451\,
            I => \ctrZ0Z_12\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__2448\,
            I => \ctrZ0Z_12\
        );

    \I__404\ : InMux
    port map (
            O => \N__2443\,
            I => ctr_cry_11
        );

    \I__403\ : InMux
    port map (
            O => \N__2440\,
            I => \N__2436\
        );

    \I__402\ : InMux
    port map (
            O => \N__2439\,
            I => \N__2433\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__2436\,
            I => \ctrZ0Z_13\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__2433\,
            I => \ctrZ0Z_13\
        );

    \I__399\ : InMux
    port map (
            O => \N__2428\,
            I => ctr_cry_12
        );

    \I__398\ : CascadeMux
    port map (
            O => \N__2425\,
            I => \N__2421\
        );

    \I__397\ : InMux
    port map (
            O => \N__2424\,
            I => \N__2418\
        );

    \I__396\ : InMux
    port map (
            O => \N__2421\,
            I => \N__2415\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__2418\,
            I => \ctrZ0Z_14\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__2415\,
            I => \ctrZ0Z_14\
        );

    \I__393\ : InMux
    port map (
            O => \N__2410\,
            I => ctr_cry_13
        );

    \I__392\ : InMux
    port map (
            O => \N__2407\,
            I => \N__2401\
        );

    \I__391\ : InMux
    port map (
            O => \N__2406\,
            I => \N__2398\
        );

    \I__390\ : InMux
    port map (
            O => \N__2405\,
            I => \N__2395\
        );

    \I__389\ : InMux
    port map (
            O => \N__2404\,
            I => \N__2392\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__2401\,
            I => \p_vLED33\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__2398\,
            I => \p_vLED33\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__2395\,
            I => \p_vLED33\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__2392\,
            I => \p_vLED33\
        );

    \I__384\ : CascadeMux
    port map (
            O => \N__2383\,
            I => \N_57_i_cascade_\
        );

    \I__383\ : CascadeMux
    port map (
            O => \N__2380\,
            I => \N__2377\
        );

    \I__382\ : InMux
    port map (
            O => \N__2377\,
            I => \N__2373\
        );

    \I__381\ : InMux
    port map (
            O => \N__2376\,
            I => \N__2370\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__2373\,
            I => \N_76\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__2370\,
            I => \N_76\
        );

    \I__378\ : InMux
    port map (
            O => \N__2365\,
            I => \N__2346\
        );

    \I__377\ : InMux
    port map (
            O => \N__2364\,
            I => \N__2346\
        );

    \I__376\ : InMux
    port map (
            O => \N__2363\,
            I => \N__2346\
        );

    \I__375\ : InMux
    port map (
            O => \N__2362\,
            I => \N__2346\
        );

    \I__374\ : InMux
    port map (
            O => \N__2361\,
            I => \N__2346\
        );

    \I__373\ : InMux
    port map (
            O => \N__2360\,
            I => \N__2346\
        );

    \I__372\ : CascadeMux
    port map (
            O => \N__2359\,
            I => \N__2340\
        );

    \I__371\ : LocalMux
    port map (
            O => \N__2346\,
            I => \N__2335\
        );

    \I__370\ : InMux
    port map (
            O => \N__2345\,
            I => \N__2328\
        );

    \I__369\ : InMux
    port map (
            O => \N__2344\,
            I => \N__2328\
        );

    \I__368\ : InMux
    port map (
            O => \N__2343\,
            I => \N__2328\
        );

    \I__367\ : InMux
    port map (
            O => \N__2340\,
            I => \N__2325\
        );

    \I__366\ : InMux
    port map (
            O => \N__2339\,
            I => \N__2320\
        );

    \I__365\ : InMux
    port map (
            O => \N__2338\,
            I => \N__2320\
        );

    \I__364\ : Odrv4
    port map (
            O => \N__2335\,
            I => \vIndexZ0Z_0\
        );

    \I__363\ : LocalMux
    port map (
            O => \N__2328\,
            I => \vIndexZ0Z_0\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__2325\,
            I => \vIndexZ0Z_0\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__2320\,
            I => \vIndexZ0Z_0\
        );

    \I__360\ : InMux
    port map (
            O => \N__2311\,
            I => \N__2307\
        );

    \I__359\ : InMux
    port map (
            O => \N__2310\,
            I => \N__2304\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__2307\,
            I => \N__2299\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__2304\,
            I => \N__2299\
        );

    \I__356\ : Odrv4
    port map (
            O => \N__2299\,
            I => \ctrZ0Z_0\
        );

    \I__355\ : InMux
    port map (
            O => \N__2296\,
            I => \bfn_9_7_0_\
        );

    \I__354\ : CascadeMux
    port map (
            O => \N__2293\,
            I => \N__2289\
        );

    \I__353\ : InMux
    port map (
            O => \N__2292\,
            I => \N__2286\
        );

    \I__352\ : InMux
    port map (
            O => \N__2289\,
            I => \N__2283\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__2286\,
            I => \ctrZ0Z_1\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__2283\,
            I => \ctrZ0Z_1\
        );

    \I__349\ : InMux
    port map (
            O => \N__2278\,
            I => ctr_cry_0
        );

    \I__348\ : InMux
    port map (
            O => \N__2275\,
            I => \N__2271\
        );

    \I__347\ : InMux
    port map (
            O => \N__2274\,
            I => \N__2268\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__2271\,
            I => \ctrZ0Z_2\
        );

    \I__345\ : LocalMux
    port map (
            O => \N__2268\,
            I => \ctrZ0Z_2\
        );

    \I__344\ : InMux
    port map (
            O => \N__2263\,
            I => ctr_cry_1
        );

    \I__343\ : InMux
    port map (
            O => \N__2260\,
            I => \N__2256\
        );

    \I__342\ : InMux
    port map (
            O => \N__2259\,
            I => \N__2253\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__2256\,
            I => \ctrZ0Z_3\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__2253\,
            I => \ctrZ0Z_3\
        );

    \I__339\ : InMux
    port map (
            O => \N__2248\,
            I => ctr_cry_2
        );

    \I__338\ : InMux
    port map (
            O => \N__2245\,
            I => \N__2241\
        );

    \I__337\ : InMux
    port map (
            O => \N__2244\,
            I => \N__2238\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__2241\,
            I => \ctrZ0Z_4\
        );

    \I__335\ : LocalMux
    port map (
            O => \N__2238\,
            I => \ctrZ0Z_4\
        );

    \I__334\ : InMux
    port map (
            O => \N__2233\,
            I => ctr_cry_3
        );

    \I__333\ : InMux
    port map (
            O => \N__2230\,
            I => \N__2226\
        );

    \I__332\ : InMux
    port map (
            O => \N__2229\,
            I => \N__2223\
        );

    \I__331\ : LocalMux
    port map (
            O => \N__2226\,
            I => \ctrZ0Z_5\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__2223\,
            I => \ctrZ0Z_5\
        );

    \I__329\ : InMux
    port map (
            O => \N__2218\,
            I => ctr_cry_4
        );

    \I__328\ : CascadeMux
    port map (
            O => \N__2215\,
            I => \N__2211\
        );

    \I__327\ : InMux
    port map (
            O => \N__2214\,
            I => \N__2208\
        );

    \I__326\ : InMux
    port map (
            O => \N__2211\,
            I => \N__2205\
        );

    \I__325\ : LocalMux
    port map (
            O => \N__2208\,
            I => \ctrZ0Z_6\
        );

    \I__324\ : LocalMux
    port map (
            O => \N__2205\,
            I => \ctrZ0Z_6\
        );

    \I__323\ : InMux
    port map (
            O => \N__2200\,
            I => ctr_cry_5
        );

    \I__322\ : InMux
    port map (
            O => \N__2197\,
            I => \N__2194\
        );

    \I__321\ : LocalMux
    port map (
            O => \N__2194\,
            I => \N__2191\
        );

    \I__320\ : Odrv4
    port map (
            O => \N__2191\,
            I => \p_vLED_cl_2_iZ0Z_0\
        );

    \I__319\ : InMux
    port map (
            O => \N__2188\,
            I => \N__2185\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__2185\,
            I => \N__2182\
        );

    \I__317\ : Odrv12
    port map (
            O => \N__2182\,
            I => \p_vLED_cl_9_iZ0Z_0\
        );

    \I__316\ : CEMux
    port map (
            O => \N__2179\,
            I => \N__2175\
        );

    \I__315\ : CEMux
    port map (
            O => \N__2178\,
            I => \N__2172\
        );

    \I__314\ : LocalMux
    port map (
            O => \N__2175\,
            I => \N__2169\
        );

    \I__313\ : LocalMux
    port map (
            O => \N__2172\,
            I => \N__2166\
        );

    \I__312\ : Odrv4
    port map (
            O => \N__2169\,
            I => \p_vLED37\
        );

    \I__311\ : Odrv4
    port map (
            O => \N__2166\,
            I => \p_vLED37\
        );

    \I__310\ : InMux
    port map (
            O => \N__2161\,
            I => \N__2141\
        );

    \I__309\ : InMux
    port map (
            O => \N__2160\,
            I => \N__2141\
        );

    \I__308\ : InMux
    port map (
            O => \N__2159\,
            I => \N__2141\
        );

    \I__307\ : InMux
    port map (
            O => \N__2158\,
            I => \N__2141\
        );

    \I__306\ : InMux
    port map (
            O => \N__2157\,
            I => \N__2141\
        );

    \I__305\ : InMux
    port map (
            O => \N__2156\,
            I => \N__2141\
        );

    \I__304\ : CascadeMux
    port map (
            O => \N__2155\,
            I => \N__2135\
        );

    \I__303\ : InMux
    port map (
            O => \N__2154\,
            I => \N__2131\
        );

    \I__302\ : LocalMux
    port map (
            O => \N__2141\,
            I => \N__2128\
        );

    \I__301\ : InMux
    port map (
            O => \N__2140\,
            I => \N__2121\
        );

    \I__300\ : InMux
    port map (
            O => \N__2139\,
            I => \N__2121\
        );

    \I__299\ : InMux
    port map (
            O => \N__2138\,
            I => \N__2121\
        );

    \I__298\ : InMux
    port map (
            O => \N__2135\,
            I => \N__2116\
        );

    \I__297\ : InMux
    port map (
            O => \N__2134\,
            I => \N__2116\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__2131\,
            I => \N__2113\
        );

    \I__295\ : Odrv4
    port map (
            O => \N__2128\,
            I => \vIndexZ0Z_2\
        );

    \I__294\ : LocalMux
    port map (
            O => \N__2121\,
            I => \vIndexZ0Z_2\
        );

    \I__293\ : LocalMux
    port map (
            O => \N__2116\,
            I => \vIndexZ0Z_2\
        );

    \I__292\ : Odrv4
    port map (
            O => \N__2113\,
            I => \vIndexZ0Z_2\
        );

    \I__291\ : CascadeMux
    port map (
            O => \N__2104\,
            I => \N__2097\
        );

    \I__290\ : CascadeMux
    port map (
            O => \N__2103\,
            I => \N__2094\
        );

    \I__289\ : CascadeMux
    port map (
            O => \N__2102\,
            I => \N__2091\
        );

    \I__288\ : CascadeMux
    port map (
            O => \N__2101\,
            I => \N__2085\
        );

    \I__287\ : CascadeMux
    port map (
            O => \N__2100\,
            I => \N__2082\
        );

    \I__286\ : InMux
    port map (
            O => \N__2097\,
            I => \N__2068\
        );

    \I__285\ : InMux
    port map (
            O => \N__2094\,
            I => \N__2068\
        );

    \I__284\ : InMux
    port map (
            O => \N__2091\,
            I => \N__2068\
        );

    \I__283\ : InMux
    port map (
            O => \N__2090\,
            I => \N__2068\
        );

    \I__282\ : InMux
    port map (
            O => \N__2089\,
            I => \N__2068\
        );

    \I__281\ : InMux
    port map (
            O => \N__2088\,
            I => \N__2068\
        );

    \I__280\ : InMux
    port map (
            O => \N__2085\,
            I => \N__2058\
        );

    \I__279\ : InMux
    port map (
            O => \N__2082\,
            I => \N__2058\
        );

    \I__278\ : InMux
    port map (
            O => \N__2081\,
            I => \N__2058\
        );

    \I__277\ : LocalMux
    port map (
            O => \N__2068\,
            I => \N__2055\
        );

    \I__276\ : InMux
    port map (
            O => \N__2067\,
            I => \N__2052\
        );

    \I__275\ : InMux
    port map (
            O => \N__2066\,
            I => \N__2049\
        );

    \I__274\ : InMux
    port map (
            O => \N__2065\,
            I => \N__2046\
        );

    \I__273\ : LocalMux
    port map (
            O => \N__2058\,
            I => \vIndexZ0Z_1\
        );

    \I__272\ : Odrv4
    port map (
            O => \N__2055\,
            I => \vIndexZ0Z_1\
        );

    \I__271\ : LocalMux
    port map (
            O => \N__2052\,
            I => \vIndexZ0Z_1\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__2049\,
            I => \vIndexZ0Z_1\
        );

    \I__269\ : LocalMux
    port map (
            O => \N__2046\,
            I => \vIndexZ0Z_1\
        );

    \I__268\ : CascadeMux
    port map (
            O => \N__2035\,
            I => \N__2027\
        );

    \I__267\ : CascadeMux
    port map (
            O => \N__2034\,
            I => \N__2024\
        );

    \I__266\ : CascadeMux
    port map (
            O => \N__2033\,
            I => \N__2021\
        );

    \I__265\ : InMux
    port map (
            O => \N__2032\,
            I => \N__2006\
        );

    \I__264\ : InMux
    port map (
            O => \N__2031\,
            I => \N__2006\
        );

    \I__263\ : InMux
    port map (
            O => \N__2030\,
            I => \N__2006\
        );

    \I__262\ : InMux
    port map (
            O => \N__2027\,
            I => \N__2006\
        );

    \I__261\ : InMux
    port map (
            O => \N__2024\,
            I => \N__2006\
        );

    \I__260\ : InMux
    port map (
            O => \N__2021\,
            I => \N__2006\
        );

    \I__259\ : CascadeMux
    port map (
            O => \N__2020\,
            I => \N__2001\
        );

    \I__258\ : CascadeMux
    port map (
            O => \N__2019\,
            I => \N__1996\
        );

    \I__257\ : LocalMux
    port map (
            O => \N__2006\,
            I => \N__1993\
        );

    \I__256\ : InMux
    port map (
            O => \N__2005\,
            I => \N__1986\
        );

    \I__255\ : InMux
    port map (
            O => \N__2004\,
            I => \N__1986\
        );

    \I__254\ : InMux
    port map (
            O => \N__2001\,
            I => \N__1986\
        );

    \I__253\ : InMux
    port map (
            O => \N__2000\,
            I => \N__1983\
        );

    \I__252\ : InMux
    port map (
            O => \N__1999\,
            I => \N__1980\
        );

    \I__251\ : InMux
    port map (
            O => \N__1996\,
            I => \N__1977\
        );

    \I__250\ : Odrv4
    port map (
            O => \N__1993\,
            I => \vIndexZ0Z_3\
        );

    \I__249\ : LocalMux
    port map (
            O => \N__1986\,
            I => \vIndexZ0Z_3\
        );

    \I__248\ : LocalMux
    port map (
            O => \N__1983\,
            I => \vIndexZ0Z_3\
        );

    \I__247\ : LocalMux
    port map (
            O => \N__1980\,
            I => \vIndexZ0Z_3\
        );

    \I__246\ : LocalMux
    port map (
            O => \N__1977\,
            I => \vIndexZ0Z_3\
        );

    \I__245\ : CascadeMux
    port map (
            O => \N__1966\,
            I => \N_76_cascade_\
        );

    \I__244\ : InMux
    port map (
            O => \N__1963\,
            I => \N__1960\
        );

    \I__243\ : LocalMux
    port map (
            O => \N__1960\,
            I => \N_57_i\
        );

    \I__242\ : CascadeMux
    port map (
            O => \N__1957\,
            I => \ballXVel12_10_cascade_\
        );

    \I__241\ : InMux
    port map (
            O => \N__1954\,
            I => \N__1951\
        );

    \I__240\ : LocalMux
    port map (
            O => \N__1951\,
            I => \ballXVel12_12\
        );

    \I__239\ : CascadeMux
    port map (
            O => \N__1948\,
            I => \ballXVel12_14_cascade_\
        );

    \I__238\ : InMux
    port map (
            O => \N__1945\,
            I => \N__1942\
        );

    \I__237\ : LocalMux
    port map (
            O => \N__1942\,
            I => \ballXVel12_11\
        );

    \I__236\ : CascadeMux
    port map (
            O => \N__1939\,
            I => \N__1933\
        );

    \I__235\ : CascadeMux
    port map (
            O => \N__1938\,
            I => \N__1928\
        );

    \I__234\ : CascadeMux
    port map (
            O => \N__1937\,
            I => \N__1922\
        );

    \I__233\ : InMux
    port map (
            O => \N__1936\,
            I => \N__1918\
        );

    \I__232\ : InMux
    port map (
            O => \N__1933\,
            I => \N__1913\
        );

    \I__231\ : InMux
    port map (
            O => \N__1932\,
            I => \N__1913\
        );

    \I__230\ : InMux
    port map (
            O => \N__1931\,
            I => \N__1904\
        );

    \I__229\ : InMux
    port map (
            O => \N__1928\,
            I => \N__1904\
        );

    \I__228\ : InMux
    port map (
            O => \N__1927\,
            I => \N__1904\
        );

    \I__227\ : InMux
    port map (
            O => \N__1926\,
            I => \N__1904\
        );

    \I__226\ : InMux
    port map (
            O => \N__1925\,
            I => \N__1897\
        );

    \I__225\ : InMux
    port map (
            O => \N__1922\,
            I => \N__1897\
        );

    \I__224\ : InMux
    port map (
            O => \N__1921\,
            I => \N__1897\
        );

    \I__223\ : LocalMux
    port map (
            O => \N__1918\,
            I => \ballXVel12\
        );

    \I__222\ : LocalMux
    port map (
            O => \N__1913\,
            I => \ballXVel12\
        );

    \I__221\ : LocalMux
    port map (
            O => \N__1904\,
            I => \ballXVel12\
        );

    \I__220\ : LocalMux
    port map (
            O => \N__1897\,
            I => \ballXVel12\
        );

    \I__219\ : InMux
    port map (
            O => \N__1888\,
            I => \N__1885\
        );

    \I__218\ : LocalMux
    port map (
            O => \N__1885\,
            I => \ballXVel12_13\
        );

    \I__217\ : IoInMux
    port map (
            O => \N__1882\,
            I => \N__1879\
        );

    \I__216\ : LocalMux
    port map (
            O => \N__1879\,
            I => \N__1876\
        );

    \I__215\ : Odrv12
    port map (
            O => \N__1876\,
            I => \N_430_i\
        );

    \I__214\ : IoInMux
    port map (
            O => \N__1873\,
            I => \N__1870\
        );

    \I__213\ : LocalMux
    port map (
            O => \N__1870\,
            I => \N__1867\
        );

    \I__212\ : Odrv12
    port map (
            O => \N__1867\,
            I => \N_428_i\
        );

    \I__211\ : InMux
    port map (
            O => \N__1864\,
            I => \N__1861\
        );

    \I__210\ : LocalMux
    port map (
            O => \N__1861\,
            I => \N_67_i\
        );

    \I__209\ : InMux
    port map (
            O => \N__1858\,
            I => \un1_vIndex_2_cry_0\
        );

    \I__208\ : InMux
    port map (
            O => \N__1855\,
            I => \un1_vIndex_2_cry_1\
        );

    \I__207\ : InMux
    port map (
            O => \N__1852\,
            I => \un1_vIndex_2_cry_2\
        );

    \I__206\ : InMux
    port map (
            O => \N__1849\,
            I => \N__1844\
        );

    \I__205\ : InMux
    port map (
            O => \N__1848\,
            I => \N__1839\
        );

    \I__204\ : InMux
    port map (
            O => \N__1847\,
            I => \N__1839\
        );

    \I__203\ : LocalMux
    port map (
            O => \N__1844\,
            I => \ballYZ0Z_0\
        );

    \I__202\ : LocalMux
    port map (
            O => \N__1839\,
            I => \ballYZ0Z_0\
        );

    \I__201\ : CascadeMux
    port map (
            O => \N__1834\,
            I => \N__1831\
        );

    \I__200\ : InMux
    port map (
            O => \N__1831\,
            I => \N__1826\
        );

    \I__199\ : InMux
    port map (
            O => \N__1830\,
            I => \N__1823\
        );

    \I__198\ : InMux
    port map (
            O => \N__1829\,
            I => \N__1820\
        );

    \I__197\ : LocalMux
    port map (
            O => \N__1826\,
            I => \ballYZ0Z_1\
        );

    \I__196\ : LocalMux
    port map (
            O => \N__1823\,
            I => \ballYZ0Z_1\
        );

    \I__195\ : LocalMux
    port map (
            O => \N__1820\,
            I => \ballYZ0Z_1\
        );

    \I__194\ : CascadeMux
    port map (
            O => \N__1813\,
            I => \ballYVel_s_1_0_0_cascade_\
        );

    \I__193\ : InMux
    port map (
            O => \N__1810\,
            I => \N__1803\
        );

    \I__192\ : InMux
    port map (
            O => \N__1809\,
            I => \N__1798\
        );

    \I__191\ : InMux
    port map (
            O => \N__1808\,
            I => \N__1798\
        );

    \I__190\ : InMux
    port map (
            O => \N__1807\,
            I => \N__1793\
        );

    \I__189\ : InMux
    port map (
            O => \N__1806\,
            I => \N__1793\
        );

    \I__188\ : LocalMux
    port map (
            O => \N__1803\,
            I => \ballYVelZ0Z_0\
        );

    \I__187\ : LocalMux
    port map (
            O => \N__1798\,
            I => \ballYVelZ0Z_0\
        );

    \I__186\ : LocalMux
    port map (
            O => \N__1793\,
            I => \ballYVelZ0Z_0\
        );

    \I__185\ : CascadeMux
    port map (
            O => \N__1786\,
            I => \N__1782\
        );

    \I__184\ : InMux
    port map (
            O => \N__1785\,
            I => \N__1778\
        );

    \I__183\ : InMux
    port map (
            O => \N__1782\,
            I => \N__1773\
        );

    \I__182\ : InMux
    port map (
            O => \N__1781\,
            I => \N__1773\
        );

    \I__181\ : LocalMux
    port map (
            O => \N__1778\,
            I => \ballYZ0Z_2\
        );

    \I__180\ : LocalMux
    port map (
            O => \N__1773\,
            I => \ballYZ0Z_2\
        );

    \I__179\ : CascadeMux
    port map (
            O => \N__1768\,
            I => \N__1764\
        );

    \I__178\ : CascadeMux
    port map (
            O => \N__1767\,
            I => \N__1760\
        );

    \I__177\ : InMux
    port map (
            O => \N__1764\,
            I => \N__1757\
        );

    \I__176\ : InMux
    port map (
            O => \N__1763\,
            I => \N__1752\
        );

    \I__175\ : InMux
    port map (
            O => \N__1760\,
            I => \N__1752\
        );

    \I__174\ : LocalMux
    port map (
            O => \N__1757\,
            I => \N__1747\
        );

    \I__173\ : LocalMux
    port map (
            O => \N__1752\,
            I => \N__1747\
        );

    \I__172\ : Odrv4
    port map (
            O => \N__1747\,
            I => \ballYZ0Z_3\
        );

    \I__171\ : InMux
    port map (
            O => \N__1744\,
            I => \N__1741\
        );

    \I__170\ : LocalMux
    port map (
            O => \N__1741\,
            I => \p_vLED37_NE_0\
        );

    \I__169\ : InMux
    port map (
            O => \N__1738\,
            I => \un1_ballX_3_cry_0\
        );

    \I__168\ : InMux
    port map (
            O => \N__1735\,
            I => \un1_ballX_3_cry_1\
        );

    \I__167\ : InMux
    port map (
            O => \N__1732\,
            I => \un1_ballX_3_cry_2\
        );

    \I__166\ : CascadeMux
    port map (
            O => \N__1729\,
            I => \ballXVel_s_1_0_0_cascade_\
        );

    \I__165\ : CascadeMux
    port map (
            O => \N__1726\,
            I => \N__1723\
        );

    \I__164\ : InMux
    port map (
            O => \N__1723\,
            I => \N__1720\
        );

    \I__163\ : LocalMux
    port map (
            O => \N__1720\,
            I => \ballXVel_RNIFI1J4_0Z0Z_0\
        );

    \I__162\ : InMux
    port map (
            O => \N__1717\,
            I => \N__1702\
        );

    \I__161\ : InMux
    port map (
            O => \N__1716\,
            I => \N__1702\
        );

    \I__160\ : InMux
    port map (
            O => \N__1715\,
            I => \N__1702\
        );

    \I__159\ : InMux
    port map (
            O => \N__1714\,
            I => \N__1702\
        );

    \I__158\ : InMux
    port map (
            O => \N__1713\,
            I => \N__1702\
        );

    \I__157\ : LocalMux
    port map (
            O => \N__1702\,
            I => \ballXVelZ0Z_0\
        );

    \I__156\ : CascadeMux
    port map (
            O => \N__1699\,
            I => \N__1696\
        );

    \I__155\ : InMux
    port map (
            O => \N__1696\,
            I => \N__1693\
        );

    \I__154\ : LocalMux
    port map (
            O => \N__1693\,
            I => \ballXVel_RNIFI1J4Z0Z_0\
        );

    \I__153\ : InMux
    port map (
            O => \N__1690\,
            I => \un1_ballY_4_cry_0\
        );

    \I__152\ : InMux
    port map (
            O => \N__1687\,
            I => \un1_ballY_4_cry_1\
        );

    \I__151\ : InMux
    port map (
            O => \N__1684\,
            I => \un1_ballY_4_cry_2\
        );

    \I__150\ : CascadeMux
    port map (
            O => \N__1681\,
            I => \N__1678\
        );

    \I__149\ : InMux
    port map (
            O => \N__1678\,
            I => \N__1675\
        );

    \I__148\ : LocalMux
    port map (
            O => \N__1675\,
            I => \ballYVel_RNIGOGN4_0Z0Z_0\
        );

    \I__147\ : CascadeMux
    port map (
            O => \N__1672\,
            I => \N__1669\
        );

    \I__146\ : InMux
    port map (
            O => \N__1669\,
            I => \N__1666\
        );

    \I__145\ : LocalMux
    port map (
            O => \N__1666\,
            I => \ballYVel_RNIGOGN4Z0Z_0\
        );

    \IN_MUX_bfv_9_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_7_0_\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => ctr_cry_7,
            carryinitout => \bfn_9_8_0_\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => ctr_cry_15,
            carryinitout => \bfn_9_9_0_\
        );

    \IN_MUX_bfv_7_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_6_0_\
        );

    \IN_MUX_bfv_8_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_6_0_\
        );

    \IN_MUX_bfv_7_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_7_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \ballY_0_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1849\,
            in2 => \N__1938\,
            in3 => \_gnd_net_\,
            lcout => \ballYZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_7_6_0_\,
            carryout => \un1_ballY_4_cry_0\,
            clk => \N__3171\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ballY_1_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1830\,
            in2 => \N__1672\,
            in3 => \N__1690\,
            lcout => \ballYZ0Z_1\,
            ltout => OPEN,
            carryin => \un1_ballY_4_cry_0\,
            carryout => \un1_ballY_4_cry_1\,
            clk => \N__3171\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ballY_2_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1785\,
            in2 => \N__1681\,
            in3 => \N__1687\,
            lcout => \ballYZ0Z_2\,
            ltout => OPEN,
            carryin => \un1_ballY_4_cry_1\,
            carryout => \un1_ballY_4_cry_2\,
            clk => \N__3171\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ballY_3_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000011101111000"
        )
    port map (
            in0 => \N__1810\,
            in1 => \N__1931\,
            in2 => \N__1768\,
            in3 => \N__1684\,
            lcout => \ballYZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3171\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ballYVel_RNIGOGN4_0_0_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1807\,
            in2 => \_gnd_net_\,
            in3 => \N__1927\,
            lcout => \ballYVel_RNIGOGN4_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ballYVel_RNIGOGN4_0_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1806\,
            in2 => \_gnd_net_\,
            in3 => \N__1926\,
            lcout => \ballYVel_RNIGOGN4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ballX_0_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2762\,
            in2 => \N__1937\,
            in3 => \_gnd_net_\,
            lcout => \ballXZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_7_7_0_\,
            carryout => \un1_ballX_3_cry_0\,
            clk => \N__3169\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ballX_1_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2811\,
            in2 => \N__1699\,
            in3 => \N__1738\,
            lcout => \ballXZ0Z_1\,
            ltout => OPEN,
            carryin => \un1_ballX_3_cry_0\,
            carryout => \un1_ballX_3_cry_1\,
            clk => \N__3169\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ballX_2_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2786\,
            in2 => \N__1726\,
            in3 => \N__1735\,
            lcout => \ballXZ0Z_2\,
            ltout => OPEN,
            carryin => \un1_ballX_3_cry_1\,
            carryout => \un1_ballX_3_cry_2\,
            clk => \N__3169\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ballX_3_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001010101101010"
        )
    port map (
            in0 => \N__2726\,
            in1 => \N__1717\,
            in2 => \N__1939\,
            in3 => \N__1732\,
            lcout => \ballXZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3169\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ballXVel_RNO_0_0_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001000000000"
        )
    port map (
            in0 => \N__1715\,
            in1 => \N__2810\,
            in2 => \N__2790\,
            in3 => \N__2763\,
            lcout => OPEN,
            ltout => \ballXVel_s_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ballXVel_0_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__2727\,
            in1 => \N__1716\,
            in2 => \N__1729\,
            in3 => \N__1925\,
            lcout => \ballXVelZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3169\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ballXVel_RNIFI1J4_0_0_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__1714\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1932\,
            lcout => \ballXVel_RNIFI1J4_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ballXVel_RNIFI1J4_0_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1713\,
            in2 => \_gnd_net_\,
            in3 => \N__1921\,
            lcout => \ballXVel_RNIFI1J4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ballY_RNIKQR82_1_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000010"
        )
    port map (
            in0 => \N__1744\,
            in1 => \N__1864\,
            in2 => \N__1834\,
            in3 => \N__2066\,
            lcout => \p_vLED37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ballY_RNIIR6I_0_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1963\,
            in2 => \N__2359\,
            in3 => \N__1847\,
            lcout => \N_67_i\,
            ltout => OPEN,
            carryin => \bfn_8_6_0_\,
            carryout => \un1_vIndex_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \vIndex_1_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2067\,
            in2 => \_gnd_net_\,
            in3 => \N__1858\,
            lcout => \vIndexZ0Z_1\,
            ltout => OPEN,
            carryin => \un1_vIndex_2_cry_0\,
            carryout => \un1_vIndex_2_cry_1\,
            clk => \N__3172\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \vIndex_2_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2155\,
            in3 => \N__1855\,
            lcout => \vIndexZ0Z_2\,
            ltout => OPEN,
            carryin => \un1_vIndex_2_cry_1\,
            carryout => \un1_vIndex_2_cry_2\,
            clk => \N__3172\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \vIndex_3_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000110100010"
        )
    port map (
            in0 => \N__2000\,
            in1 => \N__2406\,
            in2 => \N__2380\,
            in3 => \N__1852\,
            lcout => \vIndexZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3172\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ballYVel_RNO_0_0_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000001"
        )
    port map (
            in0 => \N__1848\,
            in1 => \N__1829\,
            in2 => \N__1786\,
            in3 => \N__1808\,
            lcout => OPEN,
            ltout => \ballYVel_s_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ballYVel_0_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__1809\,
            in1 => \N__1763\,
            in2 => \N__1813\,
            in3 => \N__1936\,
            lcout => \ballYVelZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3172\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ballY_RNIE1E41_3_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__1781\,
            in1 => \N__1999\,
            in2 => \N__1767\,
            in3 => \N__2134\,
            lcout => \p_vLED37_NE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_RNIDIAM_7_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2503\,
            in1 => \N__2517\,
            in2 => \N__2539\,
            in3 => \N__2484\,
            lcout => \ballXVel12_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_RNIM4UE_3_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2229\,
            in1 => \N__2244\,
            in2 => \N__2215\,
            in3 => \N__2259\,
            lcout => \ballXVel12_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_RNI05AM_18_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2310\,
            in1 => \N__2647\,
            in2 => \N__2293\,
            in3 => \N__2274\,
            lcout => OPEN,
            ltout => \ballXVel12_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_RNIOJLN1_15_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2671\,
            in1 => \N__2692\,
            in2 => \N__1957\,
            in3 => \N__2710\,
            lcout => OPEN,
            ltout => \ballXVel12_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_RNID5D94_3_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__1888\,
            in1 => \N__1954\,
            in2 => \N__1948\,
            in3 => \N__1945\,
            lcout => \ballXVel12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_RNIIQEC1_11_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2439\,
            in1 => \N__2454\,
            in2 => \N__2425\,
            in3 => \N__2469\,
            lcout => \ballXVel12_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p_vLED_obuft_RNO_9_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2188\,
            lcout => \N_430_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p_vLED_obuft_RNO_7_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2197\,
            lcout => \N_428_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p_vLED_cl_4_i_0_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__2157\,
            in1 => \N__2089\,
            in2 => \N__2034\,
            in3 => \N__2361\,
            lcout => \p_vLED_cl_4_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3181\,
            ce => \N__2179\,
            sr => \_gnd_net_\
        );

    \p_vLED_cl_i_0_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__2365\,
            in1 => \N__2032\,
            in2 => \N__2104\,
            in3 => \N__2161\,
            lcout => \p_vLED_cl_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3181\,
            ce => \N__2179\,
            sr => \_gnd_net_\
        );

    \p_vLED_cl_7_i_0_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__2363\,
            in1 => \N__2030\,
            in2 => \N__2102\,
            in3 => \N__2159\,
            lcout => \p_vLED_cl_7_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3181\,
            ce => \N__2179\,
            sr => \_gnd_net_\
        );

    \p_vLED_cl_2_i_0_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__2156\,
            in1 => \N__2088\,
            in2 => \N__2033\,
            in3 => \N__2360\,
            lcout => \p_vLED_cl_2_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3181\,
            ce => \N__2179\,
            sr => \_gnd_net_\
        );

    \p_vLED_cl_8_i_0_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__2364\,
            in1 => \N__2031\,
            in2 => \N__2103\,
            in3 => \N__2160\,
            lcout => \p_vLED_cl_8_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3181\,
            ce => \N__2179\,
            sr => \_gnd_net_\
        );

    \p_vLED_cl_6_i_0_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__2158\,
            in1 => \N__2090\,
            in2 => \N__2035\,
            in3 => \N__2362\,
            lcout => \p_vLED_cl_6_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3181\,
            ce => \N__2179\,
            sr => \_gnd_net_\
        );

    \p_vLED_cl_1_i_0_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__2138\,
            in1 => \N__2081\,
            in2 => \N__2020\,
            in3 => \N__2343\,
            lcout => \p_vLED_cl_1_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3177\,
            ce => \N__2178\,
            sr => \_gnd_net_\
        );

    \p_vLED_cl_9_i_0_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2405\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \p_vLED_cl_9_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3177\,
            ce => \N__2178\,
            sr => \_gnd_net_\
        );

    \p_vLED_cl_5_i_0_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__2345\,
            in1 => \N__2140\,
            in2 => \N__2101\,
            in3 => \N__2005\,
            lcout => \p_vLED_cl_5_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3177\,
            ce => \N__2178\,
            sr => \_gnd_net_\
        );

    \p_vLED_cl_3_i_0_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__2344\,
            in1 => \N__2139\,
            in2 => \N__2100\,
            in3 => \N__2004\,
            lcout => \p_vLED_cl_3_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3177\,
            ce => \N__2178\,
            sr => \_gnd_net_\
        );

    \vIndex_RNIUK6M_3_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__2154\,
            in1 => \N__2065\,
            in2 => \N__2019\,
            in3 => \N__2338\,
            lcout => \p_vLED33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \hIndex_RNI6JO41_1_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__3483\,
            in1 => \N__3248\,
            in2 => \N__3586\,
            in3 => \N__3379\,
            lcout => \N_76\,
            ltout => \N_76_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \vIndex_RNI48VQ1_3_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1966\,
            in3 => \N__2404\,
            lcout => \N_57_i\,
            ltout => \N_57_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \vIndex_0_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101000010010"
        )
    port map (
            in0 => \N__2339\,
            in1 => \N__2407\,
            in2 => \N__2383\,
            in3 => \N__2376\,
            lcout => \vIndexZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3175\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_0_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2311\,
            in2 => \_gnd_net_\,
            in3 => \N__2296\,
            lcout => \ctrZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_9_7_0_\,
            carryout => ctr_cry_0,
            clk => \N__3173\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_1_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2292\,
            in2 => \_gnd_net_\,
            in3 => \N__2278\,
            lcout => \ctrZ0Z_1\,
            ltout => OPEN,
            carryin => ctr_cry_0,
            carryout => ctr_cry_1,
            clk => \N__3173\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_2_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2275\,
            in2 => \_gnd_net_\,
            in3 => \N__2263\,
            lcout => \ctrZ0Z_2\,
            ltout => OPEN,
            carryin => ctr_cry_1,
            carryout => ctr_cry_2,
            clk => \N__3173\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_3_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2260\,
            in2 => \_gnd_net_\,
            in3 => \N__2248\,
            lcout => \ctrZ0Z_3\,
            ltout => OPEN,
            carryin => ctr_cry_2,
            carryout => ctr_cry_3,
            clk => \N__3173\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_4_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2245\,
            in2 => \_gnd_net_\,
            in3 => \N__2233\,
            lcout => \ctrZ0Z_4\,
            ltout => OPEN,
            carryin => ctr_cry_3,
            carryout => ctr_cry_4,
            clk => \N__3173\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_5_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2230\,
            in2 => \_gnd_net_\,
            in3 => \N__2218\,
            lcout => \ctrZ0Z_5\,
            ltout => OPEN,
            carryin => ctr_cry_4,
            carryout => ctr_cry_5,
            clk => \N__3173\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_6_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2214\,
            in2 => \_gnd_net_\,
            in3 => \N__2200\,
            lcout => \ctrZ0Z_6\,
            ltout => OPEN,
            carryin => ctr_cry_5,
            carryout => ctr_cry_6,
            clk => \N__3173\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_7_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2538\,
            in2 => \_gnd_net_\,
            in3 => \N__2521\,
            lcout => \ctrZ0Z_7\,
            ltout => OPEN,
            carryin => ctr_cry_6,
            carryout => ctr_cry_7,
            clk => \N__3173\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_8_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2518\,
            in2 => \_gnd_net_\,
            in3 => \N__2506\,
            lcout => \ctrZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_9_8_0_\,
            carryout => ctr_cry_8,
            clk => \N__3170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_9_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2502\,
            in2 => \_gnd_net_\,
            in3 => \N__2488\,
            lcout => \ctrZ0Z_9\,
            ltout => OPEN,
            carryin => ctr_cry_8,
            carryout => ctr_cry_9,
            clk => \N__3170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_10_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2485\,
            in2 => \_gnd_net_\,
            in3 => \N__2473\,
            lcout => \ctrZ0Z_10\,
            ltout => OPEN,
            carryin => ctr_cry_9,
            carryout => ctr_cry_10,
            clk => \N__3170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_11_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2470\,
            in2 => \_gnd_net_\,
            in3 => \N__2458\,
            lcout => \ctrZ0Z_11\,
            ltout => OPEN,
            carryin => ctr_cry_10,
            carryout => ctr_cry_11,
            clk => \N__3170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_12_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2455\,
            in2 => \_gnd_net_\,
            in3 => \N__2443\,
            lcout => \ctrZ0Z_12\,
            ltout => OPEN,
            carryin => ctr_cry_11,
            carryout => ctr_cry_12,
            clk => \N__3170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_13_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2440\,
            in2 => \_gnd_net_\,
            in3 => \N__2428\,
            lcout => \ctrZ0Z_13\,
            ltout => OPEN,
            carryin => ctr_cry_12,
            carryout => ctr_cry_13,
            clk => \N__3170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_14_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2424\,
            in2 => \_gnd_net_\,
            in3 => \N__2410\,
            lcout => \ctrZ0Z_14\,
            ltout => OPEN,
            carryin => ctr_cry_13,
            carryout => ctr_cry_14,
            clk => \N__3170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_15_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2709\,
            in2 => \_gnd_net_\,
            in3 => \N__2695\,
            lcout => \ctrZ0Z_15\,
            ltout => OPEN,
            carryin => ctr_cry_14,
            carryout => ctr_cry_15,
            clk => \N__3170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_16_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2688\,
            in2 => \_gnd_net_\,
            in3 => \N__2674\,
            lcout => \ctrZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => ctr_cry_16,
            clk => \N__3174\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_17_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2667\,
            in2 => \_gnd_net_\,
            in3 => \N__2653\,
            lcout => \ctrZ0Z_17\,
            ltout => OPEN,
            carryin => ctr_cry_16,
            carryout => ctr_cry_17,
            clk => \N__3174\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_18_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2646\,
            in2 => \_gnd_net_\,
            in3 => \N__2650\,
            lcout => \ctrZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3174\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p_hLED_obuft_RNO_6_LC_11_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2995\,
            lcout => \N_412_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p_vLED_obuft_RNO_8_LC_11_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__2620\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_429_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p_vLED_obuft_RNO_4_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2596\,
            lcout => \N_425_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p_vLED_obuft_RNO_3_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__2578\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_424_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p_vLED_obuft_RNO_1_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2560\,
            lcout => \N_422_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \hIndex_RNIJ9CI_1_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3341\,
            in2 => \_gnd_net_\,
            in3 => \N__3455\,
            lcout => \N_58\,
            ltout => \N_58_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \hIndex_0_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3239\,
            in2 => \N__2836\,
            in3 => \N__3570\,
            lcout => \hIndexZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3178\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \hIndex_1_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111101110000"
        )
    port map (
            in0 => \N__3568\,
            in1 => \N__3456\,
            in2 => \N__3402\,
            in3 => \N__3244\,
            lcout => \hIndexZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3178\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \hIndex_3_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000100010"
        )
    port map (
            in0 => \N__3240\,
            in1 => \N__2972\,
            in2 => \_gnd_net_\,
            in3 => \N__3571\,
            lcout => \hIndexZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3178\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \hIndex_2_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110001001100"
        )
    port map (
            in0 => \N__3569\,
            in1 => \N__3457\,
            in2 => \N__3403\,
            in3 => \N__3245\,
            lcout => \hIndexZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3178\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p_vLED_obuft_RNO_2_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2833\,
            lcout => \N_423_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ballX_RNICMG91_1_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__2812\,
            in1 => \N__3337\,
            in2 => \N__2791\,
            in3 => \N__3451\,
            lcout => \p_hLED52_NE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ballX_RNI38OK_0_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2764\,
            in2 => \_gnd_net_\,
            in3 => \N__3230\,
            lcout => \N_70_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ballX_RNIOC1J2_3_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000010"
        )
    port map (
            in0 => \N__2746\,
            in1 => \N__2740\,
            in2 => \N__2734\,
            in3 => \N__3572\,
            lcout => \p_hLED52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p_hLED_obuft_RNO_4_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__2914\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_410_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p_hLED_cl_6_i_0_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__3486\,
            in1 => \N__3285\,
            in2 => \N__3409\,
            in3 => \N__3576\,
            lcout => \p_hLED_cl_6_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3176\,
            ce => \N__3136\,
            sr => \_gnd_net_\
        );

    \p_hLED_cl_4_i_0_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__3485\,
            in1 => \N__3284\,
            in2 => \N__3408\,
            in3 => \N__3575\,
            lcout => \p_hLED_cl_4_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3176\,
            ce => \N__3136\,
            sr => \_gnd_net_\
        );

    \p_hLED_cl_12_i_0_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__3484\,
            in1 => \N__3283\,
            in2 => \N__3407\,
            in3 => \N__3574\,
            lcout => \p_hLED_cl_12_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3176\,
            ce => \N__3136\,
            sr => \_gnd_net_\
        );

    \p_hLED_cl_8_i_0_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__3573\,
            in1 => \N__3380\,
            in2 => \N__3292\,
            in3 => \N__3487\,
            lcout => \p_hLED_cl_8_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3176\,
            ce => \N__3136\,
            sr => \_gnd_net_\
        );

    \p_vLED_obuft_RNO_6_LC_12_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2908\,
            lcout => \N_427_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p_vLED_obuft_RNO_5_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2890\,
            lcout => \N_426_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p_hLED_obuft_RNO_8_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__2983\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_414_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p_vLED_obuft_RNO_0_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2860\,
            lcout => \N_421_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p_hLED_cl_7_i_0_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__3563\,
            in1 => \N__2974\,
            in2 => \_gnd_net_\,
            in3 => \N__3247\,
            lcout => \p_hLED_cl_7_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3179\,
            ce => \N__3131\,
            sr => \_gnd_net_\
        );

    \p_hLED_cl_i_0_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__3481\,
            in1 => \N__3242\,
            in2 => \N__3405\,
            in3 => \N__3567\,
            lcout => \p_hLED_cl_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3179\,
            ce => \N__3131\,
            sr => \_gnd_net_\
        );

    \p_hLED_cl_2_i_0_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__3564\,
            in1 => \N__3482\,
            in2 => \N__3406\,
            in3 => \N__3246\,
            lcout => \p_hLED_cl_2_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3179\,
            ce => \N__3131\,
            sr => \_gnd_net_\
        );

    \p_hLED_cl_1_i_0_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__2973\,
            in1 => \N__3243\,
            in2 => \_gnd_net_\,
            in3 => \N__3565\,
            lcout => \p_hLED_cl_1_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3179\,
            ce => \N__3131\,
            sr => \_gnd_net_\
        );

    \p_hLED_cl_14_i_0_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3480\,
            in1 => \N__3241\,
            in2 => \N__3404\,
            in3 => \N__3566\,
            lcout => \p_hLED_cl_14_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3179\,
            ce => \N__3131\,
            sr => \_gnd_net_\
        );

    \p_hLED_obuft_RNO_0_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__2959\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_406_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p_hLED_obuft_RNO_2_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2947\,
            lcout => \N_408_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p_hLED_obuft_RNO_1_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3592\,
            lcout => \N_407_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p_hLED_obuft_RNO_3_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3604\,
            lcout => \N_409_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p_hLED_cl_10_i_0_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__3488\,
            in1 => \N__3584\,
            in2 => \N__3289\,
            in3 => \N__3399\,
            lcout => \p_hLED_cl_10_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3180\,
            ce => \N__3135\,
            sr => \_gnd_net_\
        );

    \p_hLED_cl_9_i_0_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__3582\,
            in1 => \N__3493\,
            in2 => \N__3412\,
            in3 => \N__3282\,
            lcout => \p_hLED_cl_9_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3180\,
            ce => \N__3135\,
            sr => \_gnd_net_\
        );

    \p_hLED_cl_3_i_0_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__3581\,
            in1 => \N__3492\,
            in2 => \N__3411\,
            in3 => \N__3281\,
            lcout => \p_hLED_cl_3_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3180\,
            ce => \N__3135\,
            sr => \_gnd_net_\
        );

    \p_hLED_cl_11_i_0_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__3489\,
            in1 => \N__3583\,
            in2 => \N__3291\,
            in3 => \N__3401\,
            lcout => \p_hLED_cl_11_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3180\,
            ce => \N__3135\,
            sr => \_gnd_net_\
        );

    \p_hLED_cl_5_i_0_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__3490\,
            in1 => \N__3585\,
            in2 => \N__3290\,
            in3 => \N__3400\,
            lcout => \p_hLED_cl_5_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3180\,
            ce => \N__3135\,
            sr => \_gnd_net_\
        );

    \p_hLED_cl_13_i_0_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__3580\,
            in1 => \N__3491\,
            in2 => \N__3410\,
            in3 => \N__3280\,
            lcout => \p_hLED_cl_13_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3180\,
            ce => \N__3135\,
            sr => \_gnd_net_\
        );

    \p_hLED_obuft_RNO_10_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3103\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_416_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p_hLED_obuft_RNO_5_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3085\,
            lcout => \N_411_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p_hLED_obuft_RNO_11_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3721\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_417_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p_hLED_obuft_RNO_12_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3700\,
            lcout => \N_418_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p_hLED_obuft_RNO_7_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3676\,
            lcout => \N_413_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p_hLED_obuft_RNO_14_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3658\,
            lcout => \N_420_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p_hLED_obuft_RNO_9_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3637\,
            lcout => \N_415_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \p_hLED_obuft_RNO_13_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3619\,
            lcout => \N_419_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
